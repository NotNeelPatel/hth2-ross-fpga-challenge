module rom #(
	parameter  SIZE = 65536
	)(
	input wire clk_i,
	input wire cen_i,	
	input wire [15:0] addr_i,
	output wire[29:0] val1_o,
	output wire[29:0] val2_o
);
reg [29:0] array [SIZE];
reg [29:0] array2 [SIZE];
reg [29:0] val1_d1, val1_d2, val2_d1, val2_d2;

always @ * begin
	array2[0]=30'd212454818;
array2[1]=30'd234504581;
array2[2]=30'd229266819;
array2[3]=30'd231362949;
array2[4]=30'd229266819;
array2[5]=30'd231362949;
array2[6]=30'd231364996;
array2[7]=30'd228216193;
array2[8]=30'd231362949;
array2[9]=30'd231362949;
array2[10]=30'd230317442;
array2[11]=30'd229266819;
array2[12]=30'd229266819;
array2[13]=30'd231364996;
array2[14]=30'd231359873;
array2[15]=30'd231362949;
array2[16]=30'd234504581;
array2[17]=30'd231362949;
array2[18]=30'd231362949;
array2[19]=30'd231364996;
array2[20]=30'd229270912;
array2[21]=30'd231362949;
array2[22]=30'd231359873;
array2[23]=30'd230317442;
array2[24]=30'd231364996;
array2[25]=30'd229266819;
array2[26]=30'd231362949;
array2[27]=30'd231359873;
array2[28]=30'd231364996;
array2[29]=30'd231362949;
array2[30]=30'd230317442;
array2[31]=30'd231364996;
array2[32]=30'd234504581;
array2[33]=30'd231359873;
array2[34]=30'd231364996;
array2[35]=30'd231364996;
array2[36]=30'd230317442;
array2[37]=30'd231364996;
array2[38]=30'd231362949;
array2[39]=30'd231364996;
array2[40]=30'd231364996;
array2[41]=30'd230317442;
array2[42]=30'd231362949;
array2[43]=30'd231359873;
array2[44]=30'd234504581;
array2[45]=30'd230317442;
array2[46]=30'd231364996;
array2[47]=30'd231359873;
array2[48]=30'd229266819;
array2[49]=30'd229266819;
array2[50]=30'd231362949;
array2[51]=30'd231359873;
array2[52]=30'd231362949;
array2[53]=30'd230317442;
array2[54]=30'd231362949;
array2[55]=30'd231362949;
array2[56]=30'd231362949;
array2[57]=30'd229266819;
array2[58]=30'd231364996;
array2[59]=30'd231359873;
array2[60]=30'd231362949;
array2[61]=30'd229266819;
array2[62]=30'd231359873;
array2[63]=30'd231362949;
array2[64]=30'd229266819;
array2[65]=30'd230317442;
array2[66]=30'd231362949;
array2[67]=30'd231364996;
array2[68]=30'd231362949;
array2[69]=30'd234504581;
array2[70]=30'd231362949;
array2[71]=30'd231362949;
array2[72]=30'd229266819;
array2[73]=30'd229266819;
array2[74]=30'd229266819;
array2[75]=30'd231362949;
array2[76]=30'd231362949;
array2[77]=30'd231362949;
array2[78]=30'd231364996;
array2[79]=30'd231362949;
array2[80]=30'd231362949;
array2[81]=30'd231362949;
array2[82]=30'd230317442;
array2[83]=30'd229266819;
array2[84]=30'd231364996;
array2[85]=30'd231364996;
array2[86]=30'd231362949;
array2[87]=30'd234504581;
array2[88]=30'd231362949;
array2[89]=30'd229266819;
array2[90]=30'd229266819;
array2[91]=30'd229266819;
array2[92]=30'd231362949;
array2[93]=30'd231362949;
array2[94]=30'd234504581;
array2[95]=30'd234504581;
array2[96]=30'd212454818;
array2[97]=30'd234504581;
array2[98]=30'd231359873;
array2[99]=30'd231364996;
array2[100]=30'd229266819;
array2[101]=30'd229266819;
array2[102]=30'd231362949;
array2[103]=30'd234504581;
array2[104]=30'd231362949;
array2[105]=30'd231364996;
array2[106]=30'd229266819;
array2[107]=30'd231362949;
array2[108]=30'd231362949;
array2[109]=30'd234504581;
array2[110]=30'd231362949;
array2[111]=30'd231362949;
array2[112]=30'd231362949;
array2[113]=30'd231362949;
array2[114]=30'd234504581;
array2[115]=30'd228216193;
array2[116]=30'd231362949;
array2[117]=30'd234504581;
array2[118]=30'd231364996;
array2[119]=30'd231362949;
array2[120]=30'd229266819;
array2[121]=30'd229266819;
array2[122]=30'd229266819;
array2[123]=30'd231362949;
array2[124]=30'd231362949;
array2[125]=30'd231364996;
array2[126]=30'd231362949;
array2[127]=30'd231362949;
array2[128]=30'd234504581;
array2[129]=30'd231362949;
array2[130]=30'd231362949;
array2[131]=30'd229266819;
array2[132]=30'd229266819;
array2[133]=30'd230317442;
array2[134]=30'd231364996;
array2[135]=30'd231362949;
array2[136]=30'd230317442;
array2[137]=30'd234504581;
array2[138]=30'd229266819;
array2[139]=30'd229266819;
array2[140]=30'd231362949;
array2[141]=30'd229266819;
array2[142]=30'd231364996;
array2[143]=30'd231359873;
array2[144]=30'd234504581;
array2[145]=30'd231364996;
array2[146]=30'd234504581;
array2[147]=30'd231362949;
array2[148]=30'd231364996;
array2[149]=30'd230317442;
array2[150]=30'd231364996;
array2[151]=30'd231362949;
array2[152]=30'd234504581;
array2[153]=30'd231362949;
array2[154]=30'd231362949;
array2[155]=30'd231362949;
array2[156]=30'd230317442;
array2[157]=30'd231362949;
array2[158]=30'd228216193;
array2[159]=30'd229266819;
array2[160]=30'd231362949;
array2[161]=30'd231362949;
array2[162]=30'd231364996;
array2[163]=30'd231364996;
array2[164]=30'd231362949;
array2[165]=30'd231362949;
array2[166]=30'd234504581;
array2[167]=30'd231362949;
array2[168]=30'd229266819;
array2[169]=30'd231362949;
array2[170]=30'd231362949;
array2[171]=30'd231362949;
array2[172]=30'd231362949;
array2[173]=30'd231359873;
array2[174]=30'd231364996;
array2[175]=30'd234504581;
array2[176]=30'd231362949;
array2[177]=30'd231364996;
array2[178]=30'd231364996;
array2[179]=30'd230317442;
array2[180]=30'd231364996;
array2[181]=30'd231362949;
array2[182]=30'd231362949;
array2[183]=30'd231364996;
array2[184]=30'd228216193;
array2[185]=30'd231362949;
array2[186]=30'd231362949;
array2[187]=30'd229266819;
array2[188]=30'd229266819;
array2[189]=30'd231362949;
array2[190]=30'd229266819;
array2[191]=30'd231362949;
array2[192]=30'd212454818;
array2[193]=30'd234504581;
array2[194]=30'd230307208;
array2[195]=30'd229266819;
array2[196]=30'd229266819;
array2[197]=30'd230317442;
array2[198]=30'd229266819;
array2[199]=30'd231362949;
array2[200]=30'd231362949;
array2[201]=30'd231362949;
array2[202]=30'd230317442;
array2[203]=30'd229266819;
array2[204]=30'd230317442;
array2[205]=30'd231362949;
array2[206]=30'd231362949;
array2[207]=30'd231362949;
array2[208]=30'd231359873;
array2[209]=30'd231362949;
array2[210]=30'd230307208;
array2[211]=30'd228181405;
array2[212]=30'd232392085;
array2[213]=30'd227165569;
array2[214]=30'd229266819;
array2[215]=30'd228216193;
array2[216]=30'd228216193;
array2[217]=30'd231362949;
array2[218]=30'd231362949;
array2[219]=30'd229266819;
array2[220]=30'd229266819;
array2[221]=30'd231364996;
array2[222]=30'd230317442;
array2[223]=30'd229266819;
array2[224]=30'd230317442;
array2[225]=30'd230317442;
array2[226]=30'd231362949;
array2[227]=30'd231362949;
array2[228]=30'd231362949;
array2[229]=30'd231362949;
array2[230]=30'd229266819;
array2[231]=30'd229266819;
array2[232]=30'd229266819;
array2[233]=30'd231362949;
array2[234]=30'd231362949;
array2[235]=30'd231362949;
array2[236]=30'd231362949;
array2[237]=30'd231362949;
array2[238]=30'd231362949;
array2[239]=30'd231364996;
array2[240]=30'd231364996;
array2[241]=30'd231364996;
array2[242]=30'd231364996;
array2[243]=30'd231364996;
array2[244]=30'd229266819;
array2[245]=30'd229266819;
array2[246]=30'd231362949;
array2[247]=30'd231362949;
array2[248]=30'd231359873;
array2[249]=30'd231362949;
array2[250]=30'd229266819;
array2[251]=30'd230317442;
array2[252]=30'd231362949;
array2[253]=30'd234504581;
array2[254]=30'd256519562;
array2[255]=30'd236604812;
array2[256]=30'd231359873;
array2[257]=30'd231362949;
array2[258]=30'd230317442;
array2[259]=30'd231362949;
array2[260]=30'd231362949;
array2[261]=30'd230317442;
array2[262]=30'd231364996;
array2[263]=30'd231362949;
array2[264]=30'd231362949;
array2[265]=30'd234504581;
array2[266]=30'd231362949;
array2[267]=30'd231362949;
array2[268]=30'd231362949;
array2[269]=30'd231362949;
array2[270]=30'd231362949;
array2[271]=30'd231362949;
array2[272]=30'd229266819;
array2[273]=30'd231364996;
array2[274]=30'd231362949;
array2[275]=30'd231362949;
array2[276]=30'd231362949;
array2[277]=30'd229266819;
array2[278]=30'd230317442;
array2[279]=30'd231362949;
array2[280]=30'd231362949;
array2[281]=30'd234504581;
array2[282]=30'd231362949;
array2[283]=30'd234504581;
array2[284]=30'd231362949;
array2[285]=30'd231362949;
array2[286]=30'd231362949;
array2[287]=30'd230317442;
array2[288]=30'd212454818;
array2[289]=30'd234504581;
array2[290]=30'd228216193;
array2[291]=30'd229266819;
array2[292]=30'd229266819;
array2[293]=30'd230317442;
array2[294]=30'd229266819;
array2[295]=30'd229266819;
array2[296]=30'd231364996;
array2[297]=30'd231362949;
array2[298]=30'd234504581;
array2[299]=30'd231362949;
array2[300]=30'd229266819;
array2[301]=30'd230317442;
array2[302]=30'd229266819;
array2[303]=30'd231362949;
array2[304]=30'd231362949;
array2[305]=30'd231362949;
array2[306]=30'd230307208;
array2[307]=30'd295249323;
array2[308]=30'd295249323;
array2[309]=30'd295249323;
array2[310]=30'd295249323;
array2[311]=30'd248105365;
array2[312]=30'd227159434;
array2[313]=30'd227159434;
array2[314]=30'd227159434;
array2[315]=30'd227165569;
array2[316]=30'd229266819;
array2[317]=30'd231362949;
array2[318]=30'd231362949;
array2[319]=30'd231362949;
array2[320]=30'd229266819;
array2[321]=30'd229266819;
array2[322]=30'd230317442;
array2[323]=30'd230317442;
array2[324]=30'd231362949;
array2[325]=30'd234504581;
array2[326]=30'd229266819;
array2[327]=30'd231362949;
array2[328]=30'd229266819;
array2[329]=30'd229266819;
array2[330]=30'd229266819;
array2[331]=30'd231362949;
array2[332]=30'd234504581;
array2[333]=30'd234504581;
array2[334]=30'd231362949;
array2[335]=30'd231362949;
array2[336]=30'd231364996;
array2[337]=30'd377085336;
array2[338]=30'd377085336;
array2[339]=30'd234504581;
array2[340]=30'd231362949;
array2[341]=30'd231362949;
array2[342]=30'd231364996;
array2[343]=30'd231364996;
array2[344]=30'd228216193;
array2[345]=30'd231362949;
array2[346]=30'd231362949;
array2[347]=30'd229266819;
array2[348]=30'd229266819;
array2[349]=30'd338288022;
array2[350]=30'd603537847;
array2[351]=30'd338288022;
array2[352]=30'd227159434;
array2[353]=30'd229266819;
array2[354]=30'd231362949;
array2[355]=30'd231364996;
array2[356]=30'd228216193;
array2[357]=30'd230317442;
array2[358]=30'd231362949;
array2[359]=30'd228216193;
array2[360]=30'd229266819;
array2[361]=30'd231362949;
array2[362]=30'd230317442;
array2[363]=30'd229266819;
array2[364]=30'd231362949;
array2[365]=30'd231362949;
array2[366]=30'd231362949;
array2[367]=30'd234504581;
array2[368]=30'd231362949;
array2[369]=30'd231364996;
array2[370]=30'd234504581;
array2[371]=30'd231364996;
array2[372]=30'd229270912;
array2[373]=30'd229266819;
array2[374]=30'd230317442;
array2[375]=30'd231364996;
array2[376]=30'd229266819;
array2[377]=30'd231362949;
array2[378]=30'd231362949;
array2[379]=30'd229266819;
array2[380]=30'd231362949;
array2[381]=30'd229266819;
array2[382]=30'd231362949;
array2[383]=30'd229266819;
array2[384]=30'd212454818;
array2[385]=30'd234504581;
array2[386]=30'd228216193;
array2[387]=30'd229266819;
array2[388]=30'd231359873;
array2[389]=30'd229266819;
array2[390]=30'd231364996;
array2[391]=30'd228216193;
array2[392]=30'd231362949;
array2[393]=30'd231362949;
array2[394]=30'd231359873;
array2[395]=30'd231362949;
array2[396]=30'd231364996;
array2[397]=30'd229270912;
array2[398]=30'd231362949;
array2[399]=30'd234504581;
array2[400]=30'd234504581;
array2[401]=30'd231362949;
array2[402]=30'd227165569;
array2[403]=30'd295249323;
array2[404]=30'd356016571;
array2[405]=30'd359161273;
array2[406]=30'd359161273;
array2[407]=30'd364405173;
array2[408]=30'd312021416;
array2[409]=30'd295249323;
array2[410]=30'd295249323;
array2[411]=30'd227159434;
array2[412]=30'd221916546;
array2[413]=30'd227159434;
array2[414]=30'd230307208;
array2[415]=30'd228216193;
array2[416]=30'd228216193;
array2[417]=30'd229266819;
array2[418]=30'd231359873;
array2[419]=30'd231364996;
array2[420]=30'd231362949;
array2[421]=30'd231362949;
array2[422]=30'd229266819;
array2[423]=30'd231362949;
array2[424]=30'd228216193;
array2[425]=30'd231362949;
array2[426]=30'd228216193;
array2[427]=30'd231364996;
array2[428]=30'd229266819;
array2[429]=30'd234504581;
array2[430]=30'd272255371;
array2[431]=30'd377085336;
array2[432]=30'd231362949;
array2[433]=30'd338288022;
array2[434]=30'd338288022;
array2[435]=30'd230307208;
array2[436]=30'd377085336;
array2[437]=30'd272255371;
array2[438]=30'd227165569;
array2[439]=30'd229266819;
array2[440]=30'd229266819;
array2[441]=30'd229266819;
array2[442]=30'd229266819;
array2[443]=30'd231359873;
array2[444]=30'd231362949;
array2[445]=30'd425297329;
array2[446]=30'd719920570;
array2[447]=30'd425297329;
array2[448]=30'd231362949;
array2[449]=30'd231362949;
array2[450]=30'd228216193;
array2[451]=30'd229266819;
array2[452]=30'd231362949;
array2[453]=30'd230317442;
array2[454]=30'd231362949;
array2[455]=30'd234504581;
array2[456]=30'd231359873;
array2[457]=30'd231362949;
array2[458]=30'd229266819;
array2[459]=30'd230317442;
array2[460]=30'd231362949;
array2[461]=30'd231359873;
array2[462]=30'd231362949;
array2[463]=30'd231362949;
array2[464]=30'd231362949;
array2[465]=30'd231362949;
array2[466]=30'd231362949;
array2[467]=30'd231362949;
array2[468]=30'd229266819;
array2[469]=30'd231362949;
array2[470]=30'd229270912;
array2[471]=30'd230317442;
array2[472]=30'd231362949;
array2[473]=30'd231362949;
array2[474]=30'd229266819;
array2[475]=30'd231364996;
array2[476]=30'd229266819;
array2[477]=30'd231362949;
array2[478]=30'd231362949;
array2[479]=30'd231359873;
array2[480]=30'd212454818;
array2[481]=30'd234504581;
array2[482]=30'd227165569;
array2[483]=30'd228216193;
array2[484]=30'd231362949;
array2[485]=30'd229266819;
array2[486]=30'd230317442;
array2[487]=30'd231364996;
array2[488]=30'd228216193;
array2[489]=30'd231362949;
array2[490]=30'd234504581;
array2[491]=30'd229266819;
array2[492]=30'd229266819;
array2[493]=30'd229266819;
array2[494]=30'd229266819;
array2[495]=30'd231362949;
array2[496]=30'd231362949;
array2[497]=30'd230307208;
array2[498]=30'd228212100;
array2[499]=30'd265928088;
array2[500]=30'd356016571;
array2[501]=30'd356016571;
array2[502]=30'd356016571;
array2[503]=30'd364405173;
array2[504]=30'd364405173;
array2[505]=30'd364405173;
array2[506]=30'd356016571;
array2[507]=30'd339244483;
array2[508]=30'd312021416;
array2[509]=30'd295249323;
array2[510]=30'd220861839;
array2[511]=30'd220861839;
array2[512]=30'd230307208;
array2[513]=30'd228216193;
array2[514]=30'd228216193;
array2[515]=30'd230317442;
array2[516]=30'd231364996;
array2[517]=30'd231362949;
array2[518]=30'd229266819;
array2[519]=30'd230317442;
array2[520]=30'd231362949;
array2[521]=30'd231362949;
array2[522]=30'd231362949;
array2[523]=30'd231362949;
array2[524]=30'd229266819;
array2[525]=30'd229266819;
array2[526]=30'd272255371;
array2[527]=30'd338288022;
array2[528]=30'd234504581;
array2[529]=30'd234504581;
array2[530]=30'd231364996;
array2[531]=30'd229266819;
array2[532]=30'd338288022;
array2[533]=30'd272255371;
array2[534]=30'd231362949;
array2[535]=30'd229266819;
array2[536]=30'd230317442;
array2[537]=30'd231364996;
array2[538]=30'd228216193;
array2[539]=30'd231362949;
array2[540]=30'd234504581;
array2[541]=30'd272255371;
array2[542]=30'd472496545;
array2[543]=30'd256519562;
array2[544]=30'd227165569;
array2[545]=30'd234504581;
array2[546]=30'd231362949;
array2[547]=30'd228216193;
array2[548]=30'd230317442;
array2[549]=30'd231362949;
array2[550]=30'd231362949;
array2[551]=30'd229266819;
array2[552]=30'd231364996;
array2[553]=30'd231362949;
array2[554]=30'd231362949;
array2[555]=30'd231362949;
array2[556]=30'd229266819;
array2[557]=30'd229266819;
array2[558]=30'd229266819;
array2[559]=30'd231362949;
array2[560]=30'd231362949;
array2[561]=30'd234504581;
array2[562]=30'd234504581;
array2[563]=30'd231362949;
array2[564]=30'd231362949;
array2[565]=30'd231364996;
array2[566]=30'd231364996;
array2[567]=30'd230317442;
array2[568]=30'd230317442;
array2[569]=30'd229270912;
array2[570]=30'd231364996;
array2[571]=30'd230317442;
array2[572]=30'd230317442;
array2[573]=30'd230317442;
array2[574]=30'd231359873;
array2[575]=30'd231362949;
array2[576]=30'd212454818;
array2[577]=30'd234504581;
array2[578]=30'd227165569;
array2[579]=30'd228216193;
array2[580]=30'd231362949;
array2[581]=30'd230317442;
array2[582]=30'd229266819;
array2[583]=30'd230317442;
array2[584]=30'd230317442;
array2[585]=30'd228216193;
array2[586]=30'd231362949;
array2[587]=30'd231362949;
array2[588]=30'd229266819;
array2[589]=30'd229266819;
array2[590]=30'd229266819;
array2[591]=30'd231362949;
array2[592]=30'd230307208;
array2[593]=30'd179916222;
array2[594]=30'd179916222;
array2[595]=30'd207191473;
array2[596]=30'd339244483;
array2[597]=30'd339244483;
array2[598]=30'd464076202;
array2[599]=30'd364405173;
array2[600]=30'd359161273;
array2[601]=30'd364405173;
array2[602]=30'd364405173;
array2[603]=30'd364405173;
array2[604]=30'd356016571;
array2[605]=30'd356016571;
array2[606]=30'd339244483;
array2[607]=30'd312021416;
array2[608]=30'd228181405;
array2[609]=30'd210373000;
array2[610]=30'd232392085;
array2[611]=30'd231362949;
array2[612]=30'd231362949;
array2[613]=30'd230317442;
array2[614]=30'd231364996;
array2[615]=30'd230317442;
array2[616]=30'd231362949;
array2[617]=30'd229266819;
array2[618]=30'd229266819;
array2[619]=30'd231364996;
array2[620]=30'd229270912;
array2[621]=30'd377085336;
array2[622]=30'd338288022;
array2[623]=30'd227165569;
array2[624]=30'd234504581;
array2[625]=30'd228216193;
array2[626]=30'd230317442;
array2[627]=30'd229266819;
array2[628]=30'd230317442;
array2[629]=30'd377085336;
array2[630]=30'd377085336;
array2[631]=30'd231362949;
array2[632]=30'd231362949;
array2[633]=30'd377085336;
array2[634]=30'd603537847;
array2[635]=30'd603537847;
array2[636]=30'd472496545;
array2[637]=30'd338288022;
array2[638]=30'd603537847;
array2[639]=30'd338288022;
array2[640]=30'd377085336;
array2[641]=30'd603537847;
array2[642]=30'd603537847;
array2[643]=30'd377085336;
array2[644]=30'd228216193;
array2[645]=30'd231362949;
array2[646]=30'd230317442;
array2[647]=30'd231362949;
array2[648]=30'd229266819;
array2[649]=30'd231364996;
array2[650]=30'd231362949;
array2[651]=30'd231362949;
array2[652]=30'd231362949;
array2[653]=30'd230317442;
array2[654]=30'd231364996;
array2[655]=30'd234504581;
array2[656]=30'd234504581;
array2[657]=30'd234504581;
array2[658]=30'd231362949;
array2[659]=30'd234504581;
array2[660]=30'd231362949;
array2[661]=30'd231362949;
array2[662]=30'd231362949;
array2[663]=30'd231362949;
array2[664]=30'd229266819;
array2[665]=30'd231364996;
array2[666]=30'd229266819;
array2[667]=30'd231362949;
array2[668]=30'd231364996;
array2[669]=30'd231359873;
array2[670]=30'd231359873;
array2[671]=30'd231364996;
array2[672]=30'd212454818;
array2[673]=30'd231362949;
array2[674]=30'd227165569;
array2[675]=30'd228216193;
array2[676]=30'd229266819;
array2[677]=30'd230317442;
array2[678]=30'd231359873;
array2[679]=30'd229266819;
array2[680]=30'd229266819;
array2[681]=30'd231362949;
array2[682]=30'd231359873;
array2[683]=30'd231362949;
array2[684]=30'd230317442;
array2[685]=30'd231362949;
array2[686]=30'd231362949;
array2[687]=30'd234504581;
array2[688]=30'd269069720;
array2[689]=30'd483727963;
array2[690]=30'd645112409;
array2[691]=30'd450208341;
array2[692]=30'd444954173;
array2[693]=30'd444954173;
array2[694]=30'd381167075;
array2[695]=30'd381167075;
array2[696]=30'd356016571;
array2[697]=30'd359161273;
array2[698]=30'd356016571;
array2[699]=30'd359161273;
array2[700]=30'd356016571;
array2[701]=30'd356016571;
array2[702]=30'd356016571;
array2[703]=30'd356016571;
array2[704]=30'd339244483;
array2[705]=30'd339244483;
array2[706]=30'd312021416;
array2[707]=30'd228181405;
array2[708]=30'd221916546;
array2[709]=30'd228212100;
array2[710]=30'd230307208;
array2[711]=30'd234504581;
array2[712]=30'd229266819;
array2[713]=30'd231362949;
array2[714]=30'd228216193;
array2[715]=30'd231362949;
array2[716]=30'd231364996;
array2[717]=30'd338288022;
array2[718]=30'd338288022;
array2[719]=30'd227165569;
array2[720]=30'd231359873;
array2[721]=30'd229266819;
array2[722]=30'd231362949;
array2[723]=30'd229266819;
array2[724]=30'd231362949;
array2[725]=30'd338288022;
array2[726]=30'd338288022;
array2[727]=30'd227165569;
array2[728]=30'd231362949;
array2[729]=30'd338288022;
array2[730]=30'd532258209;
array2[731]=30'd532258209;
array2[732]=30'd464076202;
array2[733]=30'd304706973;
array2[734]=30'd532258209;
array2[735]=30'd338288022;
array2[736]=30'd338288022;
array2[737]=30'd532258209;
array2[738]=30'd553231776;
array2[739]=30'd338288022;
array2[740]=30'd231362949;
array2[741]=30'd231359873;
array2[742]=30'd231362949;
array2[743]=30'd229266819;
array2[744]=30'd229266819;
array2[745]=30'd231362949;
array2[746]=30'd229266819;
array2[747]=30'd231359873;
array2[748]=30'd231364996;
array2[749]=30'd229266819;
array2[750]=30'd231362949;
array2[751]=30'd231362949;
array2[752]=30'd231362949;
array2[753]=30'd231364996;
array2[754]=30'd231362949;
array2[755]=30'd228216193;
array2[756]=30'd231362949;
array2[757]=30'd231362949;
array2[758]=30'd229266819;
array2[759]=30'd229266819;
array2[760]=30'd229266819;
array2[761]=30'd231362949;
array2[762]=30'd231362949;
array2[763]=30'd231362949;
array2[764]=30'd231362949;
array2[765]=30'd231362949;
array2[766]=30'd231362949;
array2[767]=30'd231364996;
array2[768]=30'd212454818;
array2[769]=30'd228216193;
array2[770]=30'd234504581;
array2[771]=30'd229266819;
array2[772]=30'd231362949;
array2[773]=30'd229266819;
array2[774]=30'd231364996;
array2[775]=30'd229266819;
array2[776]=30'd228216193;
array2[777]=30'd231362949;
array2[778]=30'd229266819;
array2[779]=30'd230317442;
array2[780]=30'd231359873;
array2[781]=30'd231362949;
array2[782]=30'd231362949;
array2[783]=30'd231362949;
array2[784]=30'd295249323;
array2[785]=30'd538207812;
array2[786]=30'd729975381;
array2[787]=30'd708987491;
array2[788]=30'd805398138;
array2[789]=30'd764529268;
array2[790]=30'd538207812;
array2[791]=30'd506770009;
array2[792]=30'd389419527;
array2[793]=30'd339244483;
array2[794]=30'd339244483;
array2[795]=30'd359161273;
array2[796]=30'd356016571;
array2[797]=30'd356016571;
array2[798]=30'd356016571;
array2[799]=30'd359161273;
array2[800]=30'd364405173;
array2[801]=30'd356016571;
array2[802]=30'd356016571;
array2[803]=30'd295249323;
array2[804]=30'd232392085;
array2[805]=30'd228216193;
array2[806]=30'd231362949;
array2[807]=30'd230317442;
array2[808]=30'd231362949;
array2[809]=30'd229266819;
array2[810]=30'd231362949;
array2[811]=30'd230317442;
array2[812]=30'd231362949;
array2[813]=30'd231362949;
array2[814]=30'd272255371;
array2[815]=30'd338288022;
array2[816]=30'd231362949;
array2[817]=30'd229266819;
array2[818]=30'd230317442;
array2[819]=30'd231364996;
array2[820]=30'd338288022;
array2[821]=30'd301610387;
array2[822]=30'd231364996;
array2[823]=30'd229266819;
array2[824]=30'd229266819;
array2[825]=30'd230317442;
array2[826]=30'd229266819;
array2[827]=30'd227165569;
array2[828]=30'd231362949;
array2[829]=30'd256519562;
array2[830]=30'd472496545;
array2[831]=30'd272255371;
array2[832]=30'd227159434;
array2[833]=30'd227165569;
array2[834]=30'd231364996;
array2[835]=30'd227165569;
array2[836]=30'd231362949;
array2[837]=30'd231364996;
array2[838]=30'd231362949;
array2[839]=30'd231362949;
array2[840]=30'd231362949;
array2[841]=30'd229266819;
array2[842]=30'd231362949;
array2[843]=30'd231362949;
array2[844]=30'd231362949;
array2[845]=30'd231362949;
array2[846]=30'd231362949;
array2[847]=30'd228216193;
array2[848]=30'd230317442;
array2[849]=30'd229266819;
array2[850]=30'd231364996;
array2[851]=30'd231362949;
array2[852]=30'd231362949;
array2[853]=30'd231362949;
array2[854]=30'd230317442;
array2[855]=30'd229266819;
array2[856]=30'd229266819;
array2[857]=30'd231362949;
array2[858]=30'd229266819;
array2[859]=30'd231362949;
array2[860]=30'd234504581;
array2[861]=30'd231362949;
array2[862]=30'd231362949;
array2[863]=30'd231364996;
array2[864]=30'd212454818;
array2[865]=30'd227165569;
array2[866]=30'd231359873;
array2[867]=30'd228216193;
array2[868]=30'd230317442;
array2[869]=30'd230317442;
array2[870]=30'd229266819;
array2[871]=30'd229266819;
array2[872]=30'd231362949;
array2[873]=30'd231364996;
array2[874]=30'd231362949;
array2[875]=30'd231362949;
array2[876]=30'd234504581;
array2[877]=30'd229266819;
array2[878]=30'd229266819;
array2[879]=30'd229266819;
array2[880]=30'd257539480;
array2[881]=30'd538207812;
array2[882]=30'd729975381;
array2[883]=30'd729975381;
array2[884]=30'd790726247;
array2[885]=30'd851505800;
array2[886]=30'd851505800;
array2[887]=30'd851505800;
array2[888]=30'd646130287;
array2[889]=30'd538207812;
array2[890]=30'd506770009;
array2[891]=30'd339244483;
array2[892]=30'd339244483;
array2[893]=30'd339244483;
array2[894]=30'd356016571;
array2[895]=30'd356016571;
array2[896]=30'd359161273;
array2[897]=30'd359161273;
array2[898]=30'd356016571;
array2[899]=30'd295249323;
array2[900]=30'd227159434;
array2[901]=30'd227165569;
array2[902]=30'd229266819;
array2[903]=30'd229266819;
array2[904]=30'd231364996;
array2[905]=30'd231364996;
array2[906]=30'd231362949;
array2[907]=30'd231362949;
array2[908]=30'd231362949;
array2[909]=30'd229266819;
array2[910]=30'd301610387;
array2[911]=30'd377085336;
array2[912]=30'd231362949;
array2[913]=30'd377085336;
array2[914]=30'd377085336;
array2[915]=30'd236604812;
array2[916]=30'd377085336;
array2[917]=30'd272255371;
array2[918]=30'd231362949;
array2[919]=30'd231364996;
array2[920]=30'd231362949;
array2[921]=30'd229266819;
array2[922]=30'd231362949;
array2[923]=30'd234504581;
array2[924]=30'd229266819;
array2[925]=30'd425297329;
array2[926]=30'd719920570;
array2[927]=30'd425297329;
array2[928]=30'd231364996;
array2[929]=30'd231364996;
array2[930]=30'd231364996;
array2[931]=30'd230317442;
array2[932]=30'd231362949;
array2[933]=30'd230317442;
array2[934]=30'd231362949;
array2[935]=30'd229266819;
array2[936]=30'd229266819;
array2[937]=30'd231364996;
array2[938]=30'd231362949;
array2[939]=30'd231362949;
array2[940]=30'd234504581;
array2[941]=30'd231362949;
array2[942]=30'd229266819;
array2[943]=30'd228216193;
array2[944]=30'd231364996;
array2[945]=30'd231362949;
array2[946]=30'd231362949;
array2[947]=30'd231362949;
array2[948]=30'd231364996;
array2[949]=30'd231362949;
array2[950]=30'd231364996;
array2[951]=30'd231364996;
array2[952]=30'd231362949;
array2[953]=30'd229266819;
array2[954]=30'd231364996;
array2[955]=30'd229266819;
array2[956]=30'd231364996;
array2[957]=30'd231362949;
array2[958]=30'd228216193;
array2[959]=30'd229266819;
array2[960]=30'd212454818;
array2[961]=30'd227165569;
array2[962]=30'd231359873;
array2[963]=30'd229266819;
array2[964]=30'd231362949;
array2[965]=30'd229266819;
array2[966]=30'd229266819;
array2[967]=30'd231362949;
array2[968]=30'd231359873;
array2[969]=30'd231364996;
array2[970]=30'd231364996;
array2[971]=30'd229266819;
array2[972]=30'd231362949;
array2[973]=30'd234504581;
array2[974]=30'd231362949;
array2[975]=30'd231362949;
array2[976]=30'd220861839;
array2[977]=30'd444954173;
array2[978]=30'd737318494;
array2[979]=30'd729975381;
array2[980]=30'd737318494;
array2[981]=30'd819020415;
array2[982]=30'd858839683;
array2[983]=30'd865130113;
array2[984]=30'd858839683;
array2[985]=30'd851505800;
array2[986]=30'd819020415;
array2[987]=30'd678604396;
array2[988]=30'd646130287;
array2[989]=30'd506770009;
array2[990]=30'd281508345;
array2[991]=30'd339244483;
array2[992]=30'd356016571;
array2[993]=30'd356016571;
array2[994]=30'd339244483;
array2[995]=30'd220861839;
array2[996]=30'd228216193;
array2[997]=30'd228216193;
array2[998]=30'd231362949;
array2[999]=30'd230317442;
array2[1000]=30'd234504581;
array2[1001]=30'd229266819;
array2[1002]=30'd231364996;
array2[1003]=30'd231359873;
array2[1004]=30'd231362949;
array2[1005]=30'd231362949;
array2[1006]=30'd231359873;
array2[1007]=30'd231362949;
array2[1008]=30'd231364996;
array2[1009]=30'd377085336;
array2[1010]=30'd377085336;
array2[1011]=30'd256519562;
array2[1012]=30'd231362949;
array2[1013]=30'd231364996;
array2[1014]=30'd228216193;
array2[1015]=30'd231362949;
array2[1016]=30'd229266819;
array2[1017]=30'd231364996;
array2[1018]=30'd231362949;
array2[1019]=30'd234504581;
array2[1020]=30'd231359873;
array2[1021]=30'd338288022;
array2[1022]=30'd532258209;
array2[1023]=30'd338288022;
array2[1024]=30'd230307208;
array2[1025]=30'd229266819;
array2[1026]=30'd229266819;
array2[1027]=30'd229266819;
array2[1028]=30'd231362949;
array2[1029]=30'd231362949;
array2[1030]=30'd228216193;
array2[1031]=30'd229266819;
array2[1032]=30'd231362949;
array2[1033]=30'd231362949;
array2[1034]=30'd231362949;
array2[1035]=30'd231364996;
array2[1036]=30'd231364996;
array2[1037]=30'd231362949;
array2[1038]=30'd231362949;
array2[1039]=30'd231362949;
array2[1040]=30'd231362949;
array2[1041]=30'd231362949;
array2[1042]=30'd231362949;
array2[1043]=30'd231362949;
array2[1044]=30'd230317442;
array2[1045]=30'd231362949;
array2[1046]=30'd231362949;
array2[1047]=30'd228216193;
array2[1048]=30'd231364996;
array2[1049]=30'd231359873;
array2[1050]=30'd229266819;
array2[1051]=30'd231362949;
array2[1052]=30'd231359873;
array2[1053]=30'd231362949;
array2[1054]=30'd231362949;
array2[1055]=30'd231364996;
array2[1056]=30'd212454818;
array2[1057]=30'd234504581;
array2[1058]=30'd227165569;
array2[1059]=30'd228216193;
array2[1060]=30'd231362949;
array2[1061]=30'd230317442;
array2[1062]=30'd231359873;
array2[1063]=30'd231362949;
array2[1064]=30'd231359873;
array2[1065]=30'd229266819;
array2[1066]=30'd229266819;
array2[1067]=30'd229266819;
array2[1068]=30'd231362949;
array2[1069]=30'd231362949;
array2[1070]=30'd229266819;
array2[1071]=30'd231362949;
array2[1072]=30'd227159434;
array2[1073]=30'd444954173;
array2[1074]=30'd737318494;
array2[1075]=30'd729975381;
array2[1076]=30'd737318494;
array2[1077]=30'd819020415;
array2[1078]=30'd851505800;
array2[1079]=30'd858839683;
array2[1080]=30'd851505800;
array2[1081]=30'd851505800;
array2[1082]=30'd858839683;
array2[1083]=30'd851505800;
array2[1084]=30'd828452495;
array2[1085]=30'd764529268;
array2[1086]=30'd646130287;
array2[1087]=30'd401997362;
array2[1088]=30'd339244483;
array2[1089]=30'd359161273;
array2[1090]=30'd312021416;
array2[1091]=30'd220861839;
array2[1092]=30'd230317442;
array2[1093]=30'd229266819;
array2[1094]=30'd231364996;
array2[1095]=30'd230317442;
array2[1096]=30'd228216193;
array2[1097]=30'd231362949;
array2[1098]=30'd231362949;
array2[1099]=30'd229266819;
array2[1100]=30'd229266819;
array2[1101]=30'd229266819;
array2[1102]=30'd231362949;
array2[1103]=30'd231362949;
array2[1104]=30'd234504581;
array2[1105]=30'd234504581;
array2[1106]=30'd231364996;
array2[1107]=30'd234504581;
array2[1108]=30'd231364996;
array2[1109]=30'd231364996;
array2[1110]=30'd230317442;
array2[1111]=30'd229270912;
array2[1112]=30'd231364996;
array2[1113]=30'd230317442;
array2[1114]=30'd231364996;
array2[1115]=30'd231362949;
array2[1116]=30'd231362949;
array2[1117]=30'd231362949;
array2[1118]=30'd231359873;
array2[1119]=30'd231364996;
array2[1120]=30'd231362949;
array2[1121]=30'd231359873;
array2[1122]=30'd231362949;
array2[1123]=30'd231362949;
array2[1124]=30'd231362949;
array2[1125]=30'd231362949;
array2[1126]=30'd229266819;
array2[1127]=30'd229270912;
array2[1128]=30'd231362949;
array2[1129]=30'd234504581;
array2[1130]=30'd231362949;
array2[1131]=30'd231362949;
array2[1132]=30'd231362949;
array2[1133]=30'd229266819;
array2[1134]=30'd231362949;
array2[1135]=30'd231362949;
array2[1136]=30'd231362949;
array2[1137]=30'd234504581;
array2[1138]=30'd231362949;
array2[1139]=30'd231362949;
array2[1140]=30'd231362949;
array2[1141]=30'd231362949;
array2[1142]=30'd231362949;
array2[1143]=30'd231362949;
array2[1144]=30'd230317442;
array2[1145]=30'd231362949;
array2[1146]=30'd229266819;
array2[1147]=30'd230317442;
array2[1148]=30'd231362949;
array2[1149]=30'd231362949;
array2[1150]=30'd231362949;
array2[1151]=30'd231362949;
array2[1152]=30'd228181405;
array2[1153]=30'd227165569;
array2[1154]=30'd234504581;
array2[1155]=30'd229266819;
array2[1156]=30'd231362949;
array2[1157]=30'd230317442;
array2[1158]=30'd231362949;
array2[1159]=30'd234504581;
array2[1160]=30'd231362949;
array2[1161]=30'd231362949;
array2[1162]=30'd230317442;
array2[1163]=30'd230317442;
array2[1164]=30'd231359873;
array2[1165]=30'd231362949;
array2[1166]=30'd231362949;
array2[1167]=30'd228216193;
array2[1168]=30'd227159434;
array2[1169]=30'd444954173;
array2[1170]=30'd729975381;
array2[1171]=30'd729975381;
array2[1172]=30'd729975381;
array2[1173]=30'd737318494;
array2[1174]=30'd727851632;
array2[1175]=30'd727851632;
array2[1176]=30'd727851632;
array2[1177]=30'd727851632;
array2[1178]=30'd749877860;
array2[1179]=30'd727851632;
array2[1180]=30'd727851632;
array2[1181]=30'd727851632;
array2[1182]=30'd708987491;
array2[1183]=30'd347490866;
array2[1184]=30'd339244483;
array2[1185]=30'd339244483;
array2[1186]=30'd248105365;
array2[1187]=30'd228216193;
array2[1188]=30'd230317442;
array2[1189]=30'd231364996;
array2[1190]=30'd230317442;
array2[1191]=30'd231364996;
array2[1192]=30'd231362949;
array2[1193]=30'd229266819;
array2[1194]=30'd230317442;
array2[1195]=30'd229266819;
array2[1196]=30'd229266819;
array2[1197]=30'd231364996;
array2[1198]=30'd231362949;
array2[1199]=30'd228216193;
array2[1200]=30'd234504581;
array2[1201]=30'd231362949;
array2[1202]=30'd231362949;
array2[1203]=30'd231364996;
array2[1204]=30'd230317442;
array2[1205]=30'd231362949;
array2[1206]=30'd231364996;
array2[1207]=30'd227165569;
array2[1208]=30'd179916222;
array2[1209]=30'd150539724;
array2[1210]=30'd150539724;
array2[1211]=30'd150539724;
array2[1212]=30'd193577377;
array2[1213]=30'd232392085;
array2[1214]=30'd227159434;
array2[1215]=30'd228216193;
array2[1216]=30'd227159434;
array2[1217]=30'd228216193;
array2[1218]=30'd231364996;
array2[1219]=30'd229266819;
array2[1220]=30'd231364996;
array2[1221]=30'd229266819;
array2[1222]=30'd231362949;
array2[1223]=30'd231362949;
array2[1224]=30'd229266819;
array2[1225]=30'd231362949;
array2[1226]=30'd231362949;
array2[1227]=30'd229266819;
array2[1228]=30'd231362949;
array2[1229]=30'd231362949;
array2[1230]=30'd231362949;
array2[1231]=30'd231362949;
array2[1232]=30'd231362949;
array2[1233]=30'd231362949;
array2[1234]=30'd231364996;
array2[1235]=30'd229266819;
array2[1236]=30'd230317442;
array2[1237]=30'd229270912;
array2[1238]=30'd231362949;
array2[1239]=30'd231364996;
array2[1240]=30'd231364996;
array2[1241]=30'd229266819;
array2[1242]=30'd231362949;
array2[1243]=30'd231362949;
array2[1244]=30'd229266819;
array2[1245]=30'd231364996;
array2[1246]=30'd231362949;
array2[1247]=30'd228216193;
array2[1248]=30'd228181405;
array2[1249]=30'd227165569;
array2[1250]=30'd231362949;
array2[1251]=30'd229266819;
array2[1252]=30'd231364996;
array2[1253]=30'd231364996;
array2[1254]=30'd229266819;
array2[1255]=30'd231362949;
array2[1256]=30'd231362949;
array2[1257]=30'd231362949;
array2[1258]=30'd231362949;
array2[1259]=30'd231364996;
array2[1260]=30'd231364996;
array2[1261]=30'd231362949;
array2[1262]=30'd231359873;
array2[1263]=30'd231362949;
array2[1264]=30'd227159434;
array2[1265]=30'd383147560;
array2[1266]=30'd678604396;
array2[1267]=30'd729975381;
array2[1268]=30'd729975381;
array2[1269]=30'd729975381;
array2[1270]=30'd729975381;
array2[1271]=30'd729975381;
array2[1272]=30'd729975381;
array2[1273]=30'd737318494;
array2[1274]=30'd729975381;
array2[1275]=30'd729975381;
array2[1276]=30'd729975381;
array2[1277]=30'd737318494;
array2[1278]=30'd646130287;
array2[1279]=30'd319215128;
array2[1280]=30'd339244483;
array2[1281]=30'd339244483;
array2[1282]=30'd228181405;
array2[1283]=30'd228181405;
array2[1284]=30'd210373000;
array2[1285]=30'd248105365;
array2[1286]=30'd213516691;
array2[1287]=30'd213516691;
array2[1288]=30'd220861839;
array2[1289]=30'd228216193;
array2[1290]=30'd229266819;
array2[1291]=30'd231364996;
array2[1292]=30'd231359873;
array2[1293]=30'd231362949;
array2[1294]=30'd229266819;
array2[1295]=30'd231362949;
array2[1296]=30'd231362949;
array2[1297]=30'd231362949;
array2[1298]=30'd231364996;
array2[1299]=30'd231362949;
array2[1300]=30'd231362949;
array2[1301]=30'd234504581;
array2[1302]=30'd220861839;
array2[1303]=30'd221916546;
array2[1304]=30'd179916222;
array2[1305]=30'd150539724;
array2[1306]=30'd190356956;
array2[1307]=30'd190356956;
array2[1308]=30'd190356956;
array2[1309]=30'd190356956;
array2[1310]=30'd190356956;
array2[1311]=30'd190356956;
array2[1312]=30'd190356956;
array2[1313]=30'd212454818;
array2[1314]=30'd227159434;
array2[1315]=30'd232392085;
array2[1316]=30'd231362949;
array2[1317]=30'd227165569;
array2[1318]=30'd229266819;
array2[1319]=30'd229266819;
array2[1320]=30'd231364996;
array2[1321]=30'd229266819;
array2[1322]=30'd229266819;
array2[1323]=30'd231362949;
array2[1324]=30'd231362949;
array2[1325]=30'd231362949;
array2[1326]=30'd231364996;
array2[1327]=30'd231364996;
array2[1328]=30'd231362949;
array2[1329]=30'd231362949;
array2[1330]=30'd231362949;
array2[1331]=30'd231362949;
array2[1332]=30'd231362949;
array2[1333]=30'd231362949;
array2[1334]=30'd234504581;
array2[1335]=30'd231362949;
array2[1336]=30'd234504581;
array2[1337]=30'd231362949;
array2[1338]=30'd231364996;
array2[1339]=30'd229266819;
array2[1340]=30'd229266819;
array2[1341]=30'd231364996;
array2[1342]=30'd231359873;
array2[1343]=30'd231364996;
array2[1344]=30'd212454818;
array2[1345]=30'd231362949;
array2[1346]=30'd231362949;
array2[1347]=30'd229266819;
array2[1348]=30'd231364996;
array2[1349]=30'd230317442;
array2[1350]=30'd231364996;
array2[1351]=30'd230317442;
array2[1352]=30'd229266819;
array2[1353]=30'd230317442;
array2[1354]=30'd229266819;
array2[1355]=30'd230317442;
array2[1356]=30'd229266819;
array2[1357]=30'd231362949;
array2[1358]=30'd231362949;
array2[1359]=30'd231362949;
array2[1360]=30'd231362949;
array2[1361]=30'd207191473;
array2[1362]=30'd483727963;
array2[1363]=30'd729975381;
array2[1364]=30'd729975381;
array2[1365]=30'd729975381;
array2[1366]=30'd737318494;
array2[1367]=30'd737318494;
array2[1368]=30'd729975381;
array2[1369]=30'd729975381;
array2[1370]=30'd729975381;
array2[1371]=30'd737318494;
array2[1372]=30'd729975381;
array2[1373]=30'd708987491;
array2[1374]=30'd450208341;
array2[1375]=30'd207191473;
array2[1376]=30'd339244483;
array2[1377]=30'd359161273;
array2[1378]=30'd364405173;
array2[1379]=30'd364405173;
array2[1380]=30'd356016571;
array2[1381]=30'd356016571;
array2[1382]=30'd312021416;
array2[1383]=30'd232392085;
array2[1384]=30'd228216193;
array2[1385]=30'd228212100;
array2[1386]=30'd229270912;
array2[1387]=30'd230317442;
array2[1388]=30'd228216193;
array2[1389]=30'd231362949;
array2[1390]=30'd231362949;
array2[1391]=30'd231362949;
array2[1392]=30'd229266819;
array2[1393]=30'd229266819;
array2[1394]=30'd231362949;
array2[1395]=30'd229266819;
array2[1396]=30'd232392085;
array2[1397]=30'd195647926;
array2[1398]=30'd150539724;
array2[1399]=30'd150539724;
array2[1400]=30'd150539724;
array2[1401]=30'd249001484;
array2[1402]=30'd483727963;
array2[1403]=30'd483727963;
array2[1404]=30'd383147560;
array2[1405]=30'd407216718;
array2[1406]=30'd483727963;
array2[1407]=30'd481587821;
array2[1408]=30'd449120871;
array2[1409]=30'd383147560;
array2[1410]=30'd299264555;
array2[1411]=30'd319215128;
array2[1412]=30'd212454818;
array2[1413]=30'd213516691;
array2[1414]=30'd228216193;
array2[1415]=30'd229266819;
array2[1416]=30'd230317442;
array2[1417]=30'd231359873;
array2[1418]=30'd229266819;
array2[1419]=30'd229266819;
array2[1420]=30'd231362949;
array2[1421]=30'd231362949;
array2[1422]=30'd231362949;
array2[1423]=30'd231364996;
array2[1424]=30'd231362949;
array2[1425]=30'd231362949;
array2[1426]=30'd231359873;
array2[1427]=30'd231362949;
array2[1428]=30'd231362949;
array2[1429]=30'd231362949;
array2[1430]=30'd231362949;
array2[1431]=30'd231362949;
array2[1432]=30'd231364996;
array2[1433]=30'd234504581;
array2[1434]=30'd231362949;
array2[1435]=30'd229266819;
array2[1436]=30'd230317442;
array2[1437]=30'd231364996;
array2[1438]=30'd231362949;
array2[1439]=30'd231362949;
array2[1440]=30'd212454818;
array2[1441]=30'd234504581;
array2[1442]=30'd227165569;
array2[1443]=30'd228216193;
array2[1444]=30'd231362949;
array2[1445]=30'd230317442;
array2[1446]=30'd229266819;
array2[1447]=30'd231362949;
array2[1448]=30'd231359873;
array2[1449]=30'd230317442;
array2[1450]=30'd229266819;
array2[1451]=30'd229266819;
array2[1452]=30'd231364996;
array2[1453]=30'd231362949;
array2[1454]=30'd231362949;
array2[1455]=30'd234504581;
array2[1456]=30'd229266819;
array2[1457]=30'd193577377;
array2[1458]=30'd383147560;
array2[1459]=30'd538207812;
array2[1460]=30'd538207812;
array2[1461]=30'd538207812;
array2[1462]=30'd538207812;
array2[1463]=30'd538207812;
array2[1464]=30'd538207812;
array2[1465]=30'd538207812;
array2[1466]=30'd538207812;
array2[1467]=30'd538207812;
array2[1468]=30'd729975381;
array2[1469]=30'd645112409;
array2[1470]=30'd347490866;
array2[1471]=30'd339244483;
array2[1472]=30'd364405173;
array2[1473]=30'd356016571;
array2[1474]=30'd312021416;
array2[1475]=30'd312021416;
array2[1476]=30'd339244483;
array2[1477]=30'd356016571;
array2[1478]=30'd228181405;
array2[1479]=30'd231362949;
array2[1480]=30'd230317442;
array2[1481]=30'd228216193;
array2[1482]=30'd229270912;
array2[1483]=30'd231362949;
array2[1484]=30'd228216193;
array2[1485]=30'd231362949;
array2[1486]=30'd231362949;
array2[1487]=30'd230317442;
array2[1488]=30'd228216193;
array2[1489]=30'd231362949;
array2[1490]=30'd229266819;
array2[1491]=30'd231362949;
array2[1492]=30'd232392085;
array2[1493]=30'd179916222;
array2[1494]=30'd150539724;
array2[1495]=30'd150539724;
array2[1496]=30'd150539724;
array2[1497]=30'd249001484;
array2[1498]=30'd566515308;
array2[1499]=30'd678604396;
array2[1500]=30'd645112409;
array2[1501]=30'd538207812;
array2[1502]=30'd538207812;
array2[1503]=30'd538207812;
array2[1504]=30'd506770009;
array2[1505]=30'd481587821;
array2[1506]=30'd481587821;
array2[1507]=30'd450208341;
array2[1508]=30'd347490866;
array2[1509]=30'd281508345;
array2[1510]=30'd212454818;
array2[1511]=30'd213516691;
array2[1512]=30'd228216193;
array2[1513]=30'd231362949;
array2[1514]=30'd228216193;
array2[1515]=30'd231362949;
array2[1516]=30'd231362949;
array2[1517]=30'd231364996;
array2[1518]=30'd231362949;
array2[1519]=30'd231359873;
array2[1520]=30'd230317442;
array2[1521]=30'd231362949;
array2[1522]=30'd231362949;
array2[1523]=30'd231362949;
array2[1524]=30'd229266819;
array2[1525]=30'd229266819;
array2[1526]=30'd231364996;
array2[1527]=30'd231362949;
array2[1528]=30'd231362949;
array2[1529]=30'd231362949;
array2[1530]=30'd229266819;
array2[1531]=30'd229266819;
array2[1532]=30'd230317442;
array2[1533]=30'd229266819;
array2[1534]=30'd228216193;
array2[1535]=30'd231362949;
array2[1536]=30'd212454818;
array2[1537]=30'd234504581;
array2[1538]=30'd227165569;
array2[1539]=30'd228216193;
array2[1540]=30'd231362949;
array2[1541]=30'd230317442;
array2[1542]=30'd229266819;
array2[1543]=30'd231362949;
array2[1544]=30'd231362949;
array2[1545]=30'd229266819;
array2[1546]=30'd231362949;
array2[1547]=30'd229266819;
array2[1548]=30'd230317442;
array2[1549]=30'd231359873;
array2[1550]=30'd230317442;
array2[1551]=30'd230317442;
array2[1552]=30'd234504581;
array2[1553]=30'd213516691;
array2[1554]=30'd207191473;
array2[1555]=30'd193577377;
array2[1556]=30'd193577377;
array2[1557]=30'd193577377;
array2[1558]=30'd193577377;
array2[1559]=30'd193577377;
array2[1560]=30'd186252693;
array2[1561]=30'd193577377;
array2[1562]=30'd207191473;
array2[1563]=30'd249001484;
array2[1564]=30'd729975381;
array2[1565]=30'd538207812;
array2[1566]=30'd150539724;
array2[1567]=30'd254365107;
array2[1568]=30'd295249323;
array2[1569]=30'd254365107;
array2[1570]=30'd220861839;
array2[1571]=30'd221916546;
array2[1572]=30'd295249323;
array2[1573]=30'd295249323;
array2[1574]=30'd248105365;
array2[1575]=30'd221916546;
array2[1576]=30'd228216193;
array2[1577]=30'd229266819;
array2[1578]=30'd231364996;
array2[1579]=30'd230317442;
array2[1580]=30'd231362949;
array2[1581]=30'd234504581;
array2[1582]=30'd229266819;
array2[1583]=30'd229266819;
array2[1584]=30'd229266819;
array2[1585]=30'd230317442;
array2[1586]=30'd229266819;
array2[1587]=30'd228216193;
array2[1588]=30'd231359873;
array2[1589]=30'd232392085;
array2[1590]=30'd186252693;
array2[1591]=30'd150539724;
array2[1592]=30'd150539724;
array2[1593]=30'd150539724;
array2[1594]=30'd407216718;
array2[1595]=30'd678604396;
array2[1596]=30'd678604396;
array2[1597]=30'd729975381;
array2[1598]=30'd737318494;
array2[1599]=30'd729975381;
array2[1600]=30'd729975381;
array2[1601]=30'd645112409;
array2[1602]=30'd538207812;
array2[1603]=30'd566515308;
array2[1604]=30'd449120871;
array2[1605]=30'd407216718;
array2[1606]=30'd347490866;
array2[1607]=30'd281508345;
array2[1608]=30'd207191473;
array2[1609]=30'd207191473;
array2[1610]=30'd256519562;
array2[1611]=30'd256519562;
array2[1612]=30'd227165569;
array2[1613]=30'd229266819;
array2[1614]=30'd231362949;
array2[1615]=30'd229266819;
array2[1616]=30'd228216193;
array2[1617]=30'd229266819;
array2[1618]=30'd229266819;
array2[1619]=30'd231364996;
array2[1620]=30'd229266819;
array2[1621]=30'd231362949;
array2[1622]=30'd231362949;
array2[1623]=30'd229266819;
array2[1624]=30'd231362949;
array2[1625]=30'd231362949;
array2[1626]=30'd231362949;
array2[1627]=30'd231362949;
array2[1628]=30'd231362949;
array2[1629]=30'd229266819;
array2[1630]=30'd229266819;
array2[1631]=30'd231362949;
array2[1632]=30'd212454818;
array2[1633]=30'd231362949;
array2[1634]=30'd231362949;
array2[1635]=30'd229266819;
array2[1636]=30'd231362949;
array2[1637]=30'd230317442;
array2[1638]=30'd231362949;
array2[1639]=30'd231362949;
array2[1640]=30'd229266819;
array2[1641]=30'd231362949;
array2[1642]=30'd231362949;
array2[1643]=30'd231362949;
array2[1644]=30'd231362949;
array2[1645]=30'd231362949;
array2[1646]=30'd231362949;
array2[1647]=30'd231362949;
array2[1648]=30'd228216193;
array2[1649]=30'd229266819;
array2[1650]=30'd229266819;
array2[1651]=30'd229266819;
array2[1652]=30'd230317442;
array2[1653]=30'd231362949;
array2[1654]=30'd231362949;
array2[1655]=30'd229266819;
array2[1656]=30'd231362949;
array2[1657]=30'd231364996;
array2[1658]=30'd227159434;
array2[1659]=30'd249001484;
array2[1660]=30'd729975381;
array2[1661]=30'd538207812;
array2[1662]=30'd190356956;
array2[1663]=30'd179916222;
array2[1664]=30'd190356956;
array2[1665]=30'd179916222;
array2[1666]=30'd179916222;
array2[1667]=30'd195647926;
array2[1668]=30'd228181405;
array2[1669]=30'd228181405;
array2[1670]=30'd228181405;
array2[1671]=30'd213516691;
array2[1672]=30'd220861839;
array2[1673]=30'd227159434;
array2[1674]=30'd230307208;
array2[1675]=30'd229266819;
array2[1676]=30'd231362949;
array2[1677]=30'd231364996;
array2[1678]=30'd231362949;
array2[1679]=30'd231362949;
array2[1680]=30'd234504581;
array2[1681]=30'd229266819;
array2[1682]=30'd229266819;
array2[1683]=30'd229266819;
array2[1684]=30'd231362949;
array2[1685]=30'd231362949;
array2[1686]=30'd231364996;
array2[1687]=30'd213516691;
array2[1688]=30'd193577377;
array2[1689]=30'd124307934;
array2[1690]=30'd249001484;
array2[1691]=30'd506770009;
array2[1692]=30'd631447172;
array2[1693]=30'd646130287;
array2[1694]=30'd678604396;
array2[1695]=30'd708987491;
array2[1696]=30'd708987491;
array2[1697]=30'd729975381;
array2[1698]=30'd729975381;
array2[1699]=30'd708987491;
array2[1700]=30'd645112409;
array2[1701]=30'd566515308;
array2[1702]=30'd444954173;
array2[1703]=30'd506770009;
array2[1704]=30'd645112409;
array2[1705]=30'd538207812;
array2[1706]=30'd381167075;
array2[1707]=30'd260631016;
array2[1708]=30'd179916222;
array2[1709]=30'd212454818;
array2[1710]=30'd232392085;
array2[1711]=30'd228212100;
array2[1712]=30'd231359873;
array2[1713]=30'd231362949;
array2[1714]=30'd229266819;
array2[1715]=30'd229266819;
array2[1716]=30'd229266819;
array2[1717]=30'd229266819;
array2[1718]=30'd231364996;
array2[1719]=30'd231359873;
array2[1720]=30'd231362949;
array2[1721]=30'd231362949;
array2[1722]=30'd231364996;
array2[1723]=30'd231364996;
array2[1724]=30'd231362949;
array2[1725]=30'd231362949;
array2[1726]=30'd231362949;
array2[1727]=30'd231364996;
array2[1728]=30'd212454818;
array2[1729]=30'd234504581;
array2[1730]=30'd227165569;
array2[1731]=30'd228216193;
array2[1732]=30'd231362949;
array2[1733]=30'd230317442;
array2[1734]=30'd231359873;
array2[1735]=30'd231362949;
array2[1736]=30'd231359873;
array2[1737]=30'd230317442;
array2[1738]=30'd231362949;
array2[1739]=30'd231362949;
array2[1740]=30'd229266819;
array2[1741]=30'd229266819;
array2[1742]=30'd229270912;
array2[1743]=30'd231362949;
array2[1744]=30'd231362949;
array2[1745]=30'd234504581;
array2[1746]=30'd229266819;
array2[1747]=30'd229266819;
array2[1748]=30'd229266819;
array2[1749]=30'd229266819;
array2[1750]=30'd231362949;
array2[1751]=30'd231362949;
array2[1752]=30'd234504581;
array2[1753]=30'd231362949;
array2[1754]=30'd195647926;
array2[1755]=30'd566515308;
array2[1756]=30'd729975381;
array2[1757]=30'd678604396;
array2[1758]=30'd645112409;
array2[1759]=30'd645112409;
array2[1760]=30'd645112409;
array2[1761]=30'd645112409;
array2[1762]=30'd444954173;
array2[1763]=30'd195647926;
array2[1764]=30'd228181405;
array2[1765]=30'd254365107;
array2[1766]=30'd228181405;
array2[1767]=30'd228181405;
array2[1768]=30'd228181405;
array2[1769]=30'd228181405;
array2[1770]=30'd227159434;
array2[1771]=30'd230307208;
array2[1772]=30'd228216193;
array2[1773]=30'd231362949;
array2[1774]=30'd230317442;
array2[1775]=30'd231362949;
array2[1776]=30'd228216193;
array2[1777]=30'd227165569;
array2[1778]=30'd228212100;
array2[1779]=30'd228216193;
array2[1780]=30'd231362949;
array2[1781]=30'd230317442;
array2[1782]=30'd229266819;
array2[1783]=30'd228216193;
array2[1784]=30'd232392085;
array2[1785]=30'd212454818;
array2[1786]=30'd195647926;
array2[1787]=30'd249001484;
array2[1788]=30'd319215128;
array2[1789]=30'd566515308;
array2[1790]=30'd565444213;
array2[1791]=30'd646130287;
array2[1792]=30'd646130287;
array2[1793]=30'd678604396;
array2[1794]=30'd708987491;
array2[1795]=30'd708987491;
array2[1796]=30'd729975381;
array2[1797]=30'd708987491;
array2[1798]=30'd646130287;
array2[1799]=30'd678604396;
array2[1800]=30'd729975381;
array2[1801]=30'd708987491;
array2[1802]=30'd645112409;
array2[1803]=30'd645112409;
array2[1804]=30'd645112409;
array2[1805]=30'd444954173;
array2[1806]=30'd281508345;
array2[1807]=30'd213516691;
array2[1808]=30'd238691720;
array2[1809]=30'd231362949;
array2[1810]=30'd231362949;
array2[1811]=30'd228216193;
array2[1812]=30'd231362949;
array2[1813]=30'd231364996;
array2[1814]=30'd230317442;
array2[1815]=30'd231362949;
array2[1816]=30'd234504581;
array2[1817]=30'd231362949;
array2[1818]=30'd231359873;
array2[1819]=30'd229266819;
array2[1820]=30'd231364996;
array2[1821]=30'd228216193;
array2[1822]=30'd231362949;
array2[1823]=30'd231362949;
array2[1824]=30'd212454818;
array2[1825]=30'd227165569;
array2[1826]=30'd234504581;
array2[1827]=30'd234504581;
array2[1828]=30'd229266819;
array2[1829]=30'd229266819;
array2[1830]=30'd229266819;
array2[1831]=30'd229266819;
array2[1832]=30'd231359873;
array2[1833]=30'd229266819;
array2[1834]=30'd229266819;
array2[1835]=30'd231364996;
array2[1836]=30'd229266819;
array2[1837]=30'd231362949;
array2[1838]=30'd231364996;
array2[1839]=30'd230317442;
array2[1840]=30'd231362949;
array2[1841]=30'd229266819;
array2[1842]=30'd231362949;
array2[1843]=30'd230317442;
array2[1844]=30'd229266819;
array2[1845]=30'd231362949;
array2[1846]=30'd231362949;
array2[1847]=30'd231362949;
array2[1848]=30'd229266819;
array2[1849]=30'd231362949;
array2[1850]=30'd150539724;
array2[1851]=30'd678604396;
array2[1852]=30'd729975381;
array2[1853]=30'd729975381;
array2[1854]=30'd729975381;
array2[1855]=30'd729975381;
array2[1856]=30'd729975381;
array2[1857]=30'd645112409;
array2[1858]=30'd179916222;
array2[1859]=30'd232392085;
array2[1860]=30'd220861839;
array2[1861]=30'd228181405;
array2[1862]=30'd220861839;
array2[1863]=30'd210373000;
array2[1864]=30'd220861839;
array2[1865]=30'd248105365;
array2[1866]=30'd227159434;
array2[1867]=30'd230307208;
array2[1868]=30'd231362949;
array2[1869]=30'd229266819;
array2[1870]=30'd227165569;
array2[1871]=30'd228212100;
array2[1872]=30'd221916546;
array2[1873]=30'd228181405;
array2[1874]=30'd212454818;
array2[1875]=30'd220861839;
array2[1876]=30'd227159434;
array2[1877]=30'd227159434;
array2[1878]=30'd213516691;
array2[1879]=30'd220861839;
array2[1880]=30'd220861839;
array2[1881]=30'd220861839;
array2[1882]=30'd213516691;
array2[1883]=30'd228181405;
array2[1884]=30'd254365107;
array2[1885]=30'd281508345;
array2[1886]=30'd281508345;
array2[1887]=30'd566515308;
array2[1888]=30'd560184961;
array2[1889]=30'd560184961;
array2[1890]=30'd646130287;
array2[1891]=30'd672348794;
array2[1892]=30'd729975381;
array2[1893]=30'd729975381;
array2[1894]=30'd729975381;
array2[1895]=30'd737318494;
array2[1896]=30'd729975381;
array2[1897]=30'd737318494;
array2[1898]=30'd729975381;
array2[1899]=30'd737318494;
array2[1900]=30'd729975381;
array2[1901]=30'd678604396;
array2[1902]=30'd645112409;
array2[1903]=30'd281508345;
array2[1904]=30'd232392085;
array2[1905]=30'd227165569;
array2[1906]=30'd231364996;
array2[1907]=30'd231362949;
array2[1908]=30'd231362949;
array2[1909]=30'd231362949;
array2[1910]=30'd229266819;
array2[1911]=30'd230317442;
array2[1912]=30'd228216193;
array2[1913]=30'd231362949;
array2[1914]=30'd231362949;
array2[1915]=30'd230317442;
array2[1916]=30'd229266819;
array2[1917]=30'd231362949;
array2[1918]=30'd231362949;
array2[1919]=30'd234504581;
array2[1920]=30'd212454818;
array2[1921]=30'd234504581;
array2[1922]=30'd231362949;
array2[1923]=30'd234504581;
array2[1924]=30'd231359873;
array2[1925]=30'd229266819;
array2[1926]=30'd230317442;
array2[1927]=30'd230317442;
array2[1928]=30'd231362949;
array2[1929]=30'd231362949;
array2[1930]=30'd231362949;
array2[1931]=30'd229266819;
array2[1932]=30'd229266819;
array2[1933]=30'd230317442;
array2[1934]=30'd230317442;
array2[1935]=30'd230317442;
array2[1936]=30'd231362949;
array2[1937]=30'd229266819;
array2[1938]=30'd231364996;
array2[1939]=30'd229266819;
array2[1940]=30'd229266819;
array2[1941]=30'd229266819;
array2[1942]=30'd234504581;
array2[1943]=30'd234504581;
array2[1944]=30'd231362949;
array2[1945]=30'd230317442;
array2[1946]=30'd179916222;
array2[1947]=30'd538207812;
array2[1948]=30'd566515308;
array2[1949]=30'd645112409;
array2[1950]=30'd645112409;
array2[1951]=30'd645112409;
array2[1952]=30'd708987491;
array2[1953]=30'd566515308;
array2[1954]=30'd195647926;
array2[1955]=30'd230307208;
array2[1956]=30'd230307208;
array2[1957]=30'd232392085;
array2[1958]=30'd228216193;
array2[1959]=30'd231362949;
array2[1960]=30'd213516691;
array2[1961]=30'd232392085;
array2[1962]=30'd221916546;
array2[1963]=30'd230307208;
array2[1964]=30'd230307208;
array2[1965]=30'd230307208;
array2[1966]=30'd248105365;
array2[1967]=30'd228181405;
array2[1968]=30'd228181405;
array2[1969]=30'd254365107;
array2[1970]=30'd254365107;
array2[1971]=30'd228181405;
array2[1972]=30'd254365107;
array2[1973]=30'd254365107;
array2[1974]=30'd228181405;
array2[1975]=30'd213516691;
array2[1976]=30'd213516691;
array2[1977]=30'd220861839;
array2[1978]=30'd257539480;
array2[1979]=30'd295249323;
array2[1980]=30'd254365107;
array2[1981]=30'd260631016;
array2[1982]=30'd260631016;
array2[1983]=30'd357913199;
array2[1984]=30'd506770009;
array2[1985]=30'd483727963;
array2[1986]=30'd565444213;
array2[1987]=30'd631447172;
array2[1988]=30'd737318494;
array2[1989]=30'd729975381;
array2[1990]=30'd737318494;
array2[1991]=30'd737318494;
array2[1992]=30'd737318494;
array2[1993]=30'd729975381;
array2[1994]=30'd737318494;
array2[1995]=30'd729975381;
array2[1996]=30'd737318494;
array2[1997]=30'd737318494;
array2[1998]=30'd708987491;
array2[1999]=30'd383147560;
array2[2000]=30'd228181405;
array2[2001]=30'd228212100;
array2[2002]=30'd231364996;
array2[2003]=30'd231362949;
array2[2004]=30'd231362949;
array2[2005]=30'd229266819;
array2[2006]=30'd231359873;
array2[2007]=30'd231362949;
array2[2008]=30'd231362949;
array2[2009]=30'd231364996;
array2[2010]=30'd231364996;
array2[2011]=30'd231362949;
array2[2012]=30'd234504581;
array2[2013]=30'd234504581;
array2[2014]=30'd231362949;
array2[2015]=30'd234504581;
array2[2016]=30'd212454818;
array2[2017]=30'd228216193;
array2[2018]=30'd231364996;
array2[2019]=30'd231362949;
array2[2020]=30'd230317442;
array2[2021]=30'd231362949;
array2[2022]=30'd231364996;
array2[2023]=30'd231362949;
array2[2024]=30'd231364996;
array2[2025]=30'd231362949;
array2[2026]=30'd229266819;
array2[2027]=30'd229266819;
array2[2028]=30'd229266819;
array2[2029]=30'd230317442;
array2[2030]=30'd231364996;
array2[2031]=30'd231364996;
array2[2032]=30'd231362949;
array2[2033]=30'd231364996;
array2[2034]=30'd231362949;
array2[2035]=30'd229266819;
array2[2036]=30'd231364996;
array2[2037]=30'd230317442;
array2[2038]=30'd231364996;
array2[2039]=30'd229270912;
array2[2040]=30'd229266819;
array2[2041]=30'd229270912;
array2[2042]=30'd193577377;
array2[2043]=30'd193577377;
array2[2044]=30'd207191473;
array2[2045]=30'd212454818;
array2[2046]=30'd207191473;
array2[2047]=30'd179916222;
array2[2048]=30'd645112409;
array2[2049]=30'd444954173;
array2[2050]=30'd179916222;
array2[2051]=30'd228216193;
array2[2052]=30'd231362949;
array2[2053]=30'd231364996;
array2[2054]=30'd230317442;
array2[2055]=30'd228212100;
array2[2056]=30'd228181405;
array2[2057]=30'd228181405;
array2[2058]=30'd228181405;
array2[2059]=30'd228181405;
array2[2060]=30'd254365107;
array2[2061]=30'd295249323;
array2[2062]=30'd339244483;
array2[2063]=30'd356016571;
array2[2064]=30'd295249323;
array2[2065]=30'd254365107;
array2[2066]=30'd254365107;
array2[2067]=30'd295249323;
array2[2068]=30'd356016571;
array2[2069]=30'd356016571;
array2[2070]=30'd295249323;
array2[2071]=30'd248105365;
array2[2072]=30'd212454818;
array2[2073]=30'd195647926;
array2[2074]=30'd195647926;
array2[2075]=30'd281508345;
array2[2076]=30'd407216718;
array2[2077]=30'd518272648;
array2[2078]=30'd566515308;
array2[2079]=30'd678602388;
array2[2080]=30'd713179821;
array2[2081]=30'd713179821;
array2[2082]=30'd678602388;
array2[2083]=30'd678604396;
array2[2084]=30'd729975381;
array2[2085]=30'd729975381;
array2[2086]=30'd729975381;
array2[2087]=30'd729975381;
array2[2088]=30'd729975381;
array2[2089]=30'd737318494;
array2[2090]=30'd737318494;
array2[2091]=30'd729975381;
array2[2092]=30'd737318494;
array2[2093]=30'd737318494;
array2[2094]=30'd729975381;
array2[2095]=30'd645112409;
array2[2096]=30'd249001484;
array2[2097]=30'd227159434;
array2[2098]=30'd227165569;
array2[2099]=30'd231362949;
array2[2100]=30'd229266819;
array2[2101]=30'd229266819;
array2[2102]=30'd229266819;
array2[2103]=30'd231362949;
array2[2104]=30'd229266819;
array2[2105]=30'd231362949;
array2[2106]=30'd231364996;
array2[2107]=30'd230317442;
array2[2108]=30'd231362949;
array2[2109]=30'd231362949;
array2[2110]=30'd229266819;
array2[2111]=30'd231362949;
array2[2112]=30'd207191473;
array2[2113]=30'd240774546;
array2[2114]=30'd232392085;
array2[2115]=30'd227165569;
array2[2116]=30'd228216193;
array2[2117]=30'd230317442;
array2[2118]=30'd229266819;
array2[2119]=30'd229266819;
array2[2120]=30'd229266819;
array2[2121]=30'd230317442;
array2[2122]=30'd229266819;
array2[2123]=30'd231362949;
array2[2124]=30'd230317442;
array2[2125]=30'd229270912;
array2[2126]=30'd232392085;
array2[2127]=30'd232392085;
array2[2128]=30'd232392085;
array2[2129]=30'd232392085;
array2[2130]=30'd232392085;
array2[2131]=30'd227159434;
array2[2132]=30'd234499470;
array2[2133]=30'd234499470;
array2[2134]=30'd234499470;
array2[2135]=30'd234499470;
array2[2136]=30'd232392085;
array2[2137]=30'd232392085;
array2[2138]=30'd227165569;
array2[2139]=30'd227165569;
array2[2140]=30'd228216193;
array2[2141]=30'd231362949;
array2[2142]=30'd227165569;
array2[2143]=30'd179916222;
array2[2144]=30'd444954173;
array2[2145]=30'd190356956;
array2[2146]=30'd212454818;
array2[2147]=30'd229266819;
array2[2148]=30'd229266819;
array2[2149]=30'd227159434;
array2[2150]=30'd232392085;
array2[2151]=30'd213516691;
array2[2152]=30'd267996623;
array2[2153]=30'd254365107;
array2[2154]=30'd267996623;
array2[2155]=30'd339244483;
array2[2156]=30'd339244483;
array2[2157]=30'd381167075;
array2[2158]=30'd381167075;
array2[2159]=30'd381167075;
array2[2160]=30'd295249323;
array2[2161]=30'd295249323;
array2[2162]=30'd254365107;
array2[2163]=30'd190356956;
array2[2164]=30'd281508345;
array2[2165]=30'd281508345;
array2[2166]=30'd281508345;
array2[2167]=30'd179916222;
array2[2168]=30'd190356956;
array2[2169]=30'd375721588;
array2[2170]=30'd481587821;
array2[2171]=30'd566515308;
array2[2172]=30'd678602388;
array2[2173]=30'd770812573;
array2[2174]=30'd770812573;
array2[2175]=30'd770812573;
array2[2176]=30'd770812573;
array2[2177]=30'd805398138;
array2[2178]=30'd805398138;
array2[2179]=30'd764529268;
array2[2180]=30'd727851632;
array2[2181]=30'd737318494;
array2[2182]=30'd708987491;
array2[2183]=30'd729975381;
array2[2184]=30'd729975381;
array2[2185]=30'd737318494;
array2[2186]=30'd729975381;
array2[2187]=30'd729975381;
array2[2188]=30'd737318494;
array2[2189]=30'd737318494;
array2[2190]=30'd729975381;
array2[2191]=30'd708987491;
array2[2192]=30'd483727963;
array2[2193]=30'd193577377;
array2[2194]=30'd230307208;
array2[2195]=30'd227165569;
array2[2196]=30'd231362949;
array2[2197]=30'd229266819;
array2[2198]=30'd231362949;
array2[2199]=30'd231362949;
array2[2200]=30'd231362949;
array2[2201]=30'd228216193;
array2[2202]=30'd231359873;
array2[2203]=30'd231362949;
array2[2204]=30'd229266819;
array2[2205]=30'd229266819;
array2[2206]=30'd230317442;
array2[2207]=30'd231362949;
array2[2208]=30'd390446940;
array2[2209]=30'd461700935;
array2[2210]=30'd451191548;
array2[2211]=30'd284737060;
array2[2212]=30'd280568333;
array2[2213]=30'd280568333;
array2[2214]=30'd280568333;
array2[2215]=30'd280568333;
array2[2216]=30'd280568333;
array2[2217]=30'd280568333;
array2[2218]=30'd280568333;
array2[2219]=30'd280568333;
array2[2220]=30'd280568333;
array2[2221]=30'd302506616;
array2[2222]=30'd461700935;
array2[2223]=30'd461700935;
array2[2224]=30'd461700935;
array2[2225]=30'd461700935;
array2[2226]=30'd461700935;
array2[2227]=30'd461700935;
array2[2228]=30'd461700935;
array2[2229]=30'd461700935;
array2[2230]=30'd461700935;
array2[2231]=30'd461700935;
array2[2232]=30'd461700935;
array2[2233]=30'd390446940;
array2[2234]=30'd307771998;
array2[2235]=30'd280568333;
array2[2236]=30'd280568333;
array2[2237]=30'd280568333;
array2[2238]=30'd280568333;
array2[2239]=30'd190356956;
array2[2240]=30'd347490866;
array2[2241]=30'd265736724;
array2[2242]=30'd179916222;
array2[2243]=30'd179916222;
array2[2244]=30'd179916222;
array2[2245]=30'd287786593;
array2[2246]=30'd302506616;
array2[2247]=30'd390446940;
array2[2248]=30'd461700935;
array2[2249]=30'd390446940;
array2[2250]=30'd390446940;
array2[2251]=30'd461700935;
array2[2252]=30'd409311115;
array2[2253]=30'd461700935;
array2[2254]=30'd461700935;
array2[2255]=30'd395649781;
array2[2256]=30'd281508345;
array2[2257]=30'd190356956;
array2[2258]=30'd249001484;
array2[2259]=30'd518272648;
array2[2260]=30'd631447172;
array2[2261]=30'd566515308;
array2[2262]=30'd357913199;
array2[2263]=30'd295074390;
array2[2264]=30'd338018898;
array2[2265]=30'd631447172;
array2[2266]=30'd677571193;
array2[2267]=30'd764529268;
array2[2268]=30'd828452495;
array2[2269]=30'd828452495;
array2[2270]=30'd851505800;
array2[2271]=30'd851505800;
array2[2272]=30'd851505800;
array2[2273]=30'd851505800;
array2[2274]=30'd805398138;
array2[2275]=30'd768729747;
array2[2276]=30'd764529268;
array2[2277]=30'd764529268;
array2[2278]=30'd737318494;
array2[2279]=30'd737318494;
array2[2280]=30'd729975381;
array2[2281]=30'd737318494;
array2[2282]=30'd729975381;
array2[2283]=30'd737318494;
array2[2284]=30'd645112409;
array2[2285]=30'd401997362;
array2[2286]=30'd645112409;
array2[2287]=30'd737318494;
array2[2288]=30'd645112409;
array2[2289]=30'd195647926;
array2[2290]=30'd228216193;
array2[2291]=30'd229266819;
array2[2292]=30'd229266819;
array2[2293]=30'd229266819;
array2[2294]=30'd231359873;
array2[2295]=30'd231362949;
array2[2296]=30'd231359873;
array2[2297]=30'd228216193;
array2[2298]=30'd229266819;
array2[2299]=30'd231364996;
array2[2300]=30'd231362949;
array2[2301]=30'd231362949;
array2[2302]=30'd231362949;
array2[2303]=30'd231362949;
array2[2304]=30'd409311115;
array2[2305]=30'd426044336;
array2[2306]=30'd429185963;
array2[2307]=30'd409311115;
array2[2308]=30'd409311115;
array2[2309]=30'd409311115;
array2[2310]=30'd409311115;
array2[2311]=30'd409311115;
array2[2312]=30'd409311115;
array2[2313]=30'd409311115;
array2[2314]=30'd409311115;
array2[2315]=30'd409311115;
array2[2316]=30'd409311115;
array2[2317]=30'd429185963;
array2[2318]=30'd423950257;
array2[2319]=30'd423950257;
array2[2320]=30'd423950257;
array2[2321]=30'd423950257;
array2[2322]=30'd423950257;
array2[2323]=30'd426044336;
array2[2324]=30'd423950257;
array2[2325]=30'd426044336;
array2[2326]=30'd423950257;
array2[2327]=30'd426044336;
array2[2328]=30'd423950257;
array2[2329]=30'd429185963;
array2[2330]=30'd429185963;
array2[2331]=30'd409311115;
array2[2332]=30'd409311115;
array2[2333]=30'd409311115;
array2[2334]=30'd357996288;
array2[2335]=30'd339090072;
array2[2336]=30'd380968597;
array2[2337]=30'd380968597;
array2[2338]=30'd380968597;
array2[2339]=30'd380968597;
array2[2340]=30'd380968597;
array2[2341]=30'd380968597;
array2[2342]=30'd287786593;
array2[2343]=30'd429185963;
array2[2344]=30'd423950257;
array2[2345]=30'd409311115;
array2[2346]=30'd493111164;
array2[2347]=30'd493111164;
array2[2348]=30'd461700935;
array2[2349]=30'd357913199;
array2[2350]=30'd331763301;
array2[2351]=30'd566515308;
array2[2352]=30'd727851632;
array2[2353]=30'd727851632;
array2[2354]=30'd727851632;
array2[2355]=30'd805398138;
array2[2356]=30'd828452495;
array2[2357]=30'd678602388;
array2[2358]=30'd481587821;
array2[2359]=30'd434416250;
array2[2360]=30'd434416250;
array2[2361]=30'd727851632;
array2[2362]=30'd727851632;
array2[2363]=30'd764529268;
array2[2364]=30'd851505800;
array2[2365]=30'd851505800;
array2[2366]=30'd851505800;
array2[2367]=30'd851505800;
array2[2368]=30'd858839683;
array2[2369]=30'd858839683;
array2[2370]=30'd828452495;
array2[2371]=30'd805398138;
array2[2372]=30'd805398138;
array2[2373]=30'd828452495;
array2[2374]=30'd828452495;
array2[2375]=30'd828452495;
array2[2376]=30'd764529268;
array2[2377]=30'd727851632;
array2[2378]=30'd708987491;
array2[2379]=30'd737318494;
array2[2380]=30'd566515308;
array2[2381]=30'd195647926;
array2[2382]=30'd566515308;
array2[2383]=30'd737318494;
array2[2384]=30'd645112409;
array2[2385]=30'd195647926;
array2[2386]=30'd227159434;
array2[2387]=30'd231359873;
array2[2388]=30'd230317442;
array2[2389]=30'd231362949;
array2[2390]=30'd231364996;
array2[2391]=30'd231362949;
array2[2392]=30'd231362949;
array2[2393]=30'd234504581;
array2[2394]=30'd229266819;
array2[2395]=30'd229266819;
array2[2396]=30'd229266819;
array2[2397]=30'd231362949;
array2[2398]=30'd228216193;
array2[2399]=30'd231362949;
array2[2400]=30'd461700935;
array2[2401]=30'd426044336;
array2[2402]=30'd426044336;
array2[2403]=30'd426044336;
array2[2404]=30'd426044336;
array2[2405]=30'd426044336;
array2[2406]=30'd426044336;
array2[2407]=30'd426044336;
array2[2408]=30'd426044336;
array2[2409]=30'd426044336;
array2[2410]=30'd426044336;
array2[2411]=30'd426044336;
array2[2412]=30'd426044336;
array2[2413]=30'd426044336;
array2[2414]=30'd423950257;
array2[2415]=30'd423950257;
array2[2416]=30'd426044336;
array2[2417]=30'd426044336;
array2[2418]=30'd423950257;
array2[2419]=30'd426044336;
array2[2420]=30'd426044336;
array2[2421]=30'd423950257;
array2[2422]=30'd426044336;
array2[2423]=30'd426044336;
array2[2424]=30'd423950257;
array2[2425]=30'd426044336;
array2[2426]=30'd423950257;
array2[2427]=30'd426044336;
array2[2428]=30'd426044336;
array2[2429]=30'd426044336;
array2[2430]=30'd395649781;
array2[2431]=30'd339090072;
array2[2432]=30'd380968597;
array2[2433]=30'd380968597;
array2[2434]=30'd380968597;
array2[2435]=30'd380968597;
array2[2436]=30'd380968597;
array2[2437]=30'd331763301;
array2[2438]=30'd409311115;
array2[2439]=30'd426044336;
array2[2440]=30'd409311115;
array2[2441]=30'd493111164;
array2[2442]=30'd493111164;
array2[2443]=30'd461700935;
array2[2444]=30'd375721588;
array2[2445]=30'd449120871;
array2[2446]=30'd449120871;
array2[2447]=30'd677571193;
array2[2448]=30'd770816666;
array2[2449]=30'd764529268;
array2[2450]=30'd768729747;
array2[2451]=30'd828452495;
array2[2452]=30'd858839683;
array2[2453]=30'd762499681;
array2[2454]=30'd481587821;
array2[2455]=30'd450208341;
array2[2456]=30'd434416250;
array2[2457]=30'd764529268;
array2[2458]=30'd805398138;
array2[2459]=30'd828452495;
array2[2460]=30'd805398138;
array2[2461]=30'd828452495;
array2[2462]=30'd851505800;
array2[2463]=30'd851505800;
array2[2464]=30'd851505800;
array2[2465]=30'd858839683;
array2[2466]=30'd858839683;
array2[2467]=30'd851505800;
array2[2468]=30'd828452495;
array2[2469]=30'd851505800;
array2[2470]=30'd858839683;
array2[2471]=30'd858839683;
array2[2472]=30'd858839683;
array2[2473]=30'd828452495;
array2[2474]=30'd762499681;
array2[2475]=30'd727851632;
array2[2476]=30'd566515308;
array2[2477]=30'd150539724;
array2[2478]=30'd538207812;
array2[2479]=30'd729975381;
array2[2480]=30'd645112409;
array2[2481]=30'd179916222;
array2[2482]=30'd232392085;
array2[2483]=30'd229266819;
array2[2484]=30'd228216193;
array2[2485]=30'd231364996;
array2[2486]=30'd231362949;
array2[2487]=30'd231362949;
array2[2488]=30'd227165569;
array2[2489]=30'd227165569;
array2[2490]=30'd229266819;
array2[2491]=30'd229266819;
array2[2492]=30'd230317442;
array2[2493]=30'd228216193;
array2[2494]=30'd231362949;
array2[2495]=30'd234504581;
array2[2496]=30'd646169309;
array2[2497]=30'd672324351;
array2[2498]=30'd582196031;
array2[2499]=30'd435467177;
array2[2500]=30'd435467177;
array2[2501]=30'd426044336;
array2[2502]=30'd426044336;
array2[2503]=30'd426044336;
array2[2504]=30'd426044336;
array2[2505]=30'd426044336;
array2[2506]=30'd426044336;
array2[2507]=30'd426044336;
array2[2508]=30'd426044336;
array2[2509]=30'd493111164;
array2[2510]=30'd672324351;
array2[2511]=30'd672324351;
array2[2512]=30'd672324351;
array2[2513]=30'd672324351;
array2[2514]=30'd672324351;
array2[2515]=30'd672324351;
array2[2516]=30'd672324351;
array2[2517]=30'd672324351;
array2[2518]=30'd672324351;
array2[2519]=30'd672324351;
array2[2520]=30'd672324351;
array2[2521]=30'd635645720;
array2[2522]=30'd435467177;
array2[2523]=30'd426044336;
array2[2524]=30'd426044336;
array2[2525]=30'd426044336;
array2[2526]=30'd390446940;
array2[2527]=30'd357996288;
array2[2528]=30'd357996288;
array2[2529]=30'd380968597;
array2[2530]=30'd357996288;
array2[2531]=30'd328674981;
array2[2532]=30'd380968597;
array2[2533]=30'd331763301;
array2[2534]=30'd646169309;
array2[2535]=30'd646169309;
array2[2536]=30'd672324351;
array2[2537]=30'd646169309;
array2[2538]=30'd518272648;
array2[2539]=30'd483727963;
array2[2540]=30'd434416250;
array2[2541]=30'd481587821;
array2[2542]=30'd481587821;
array2[2543]=30'd606320275;
array2[2544]=30'd770812573;
array2[2545]=30'd819020415;
array2[2546]=30'd819020415;
array2[2547]=30'd851505800;
array2[2548]=30'd858839683;
array2[2549]=30'd768729747;
array2[2550]=30'd518272648;
array2[2551]=30'd434416250;
array2[2552]=30'd434416250;
array2[2553]=30'd764529268;
array2[2554]=30'd805398138;
array2[2555]=30'd851505800;
array2[2556]=30'd828452495;
array2[2557]=30'd790726247;
array2[2558]=30'd805398138;
array2[2559]=30'd819020415;
array2[2560]=30'd828452495;
array2[2561]=30'd851505800;
array2[2562]=30'd851505800;
array2[2563]=30'd858839683;
array2[2564]=30'd858839683;
array2[2565]=30'd851505800;
array2[2566]=30'd858839683;
array2[2567]=30'd858839683;
array2[2568]=30'd858839683;
array2[2569]=30'd828452495;
array2[2570]=30'd770812573;
array2[2571]=30'd768729747;
array2[2572]=30'd565444213;
array2[2573]=30'd284737060;
array2[2574]=30'd566515308;
array2[2575]=30'd737318494;
array2[2576]=30'd646130287;
array2[2577]=30'd450208341;
array2[2578]=30'd179916222;
array2[2579]=30'd220861839;
array2[2580]=30'd229266819;
array2[2581]=30'd229266819;
array2[2582]=30'd231364996;
array2[2583]=30'd231364996;
array2[2584]=30'd231362949;
array2[2585]=30'd234504581;
array2[2586]=30'd229266819;
array2[2587]=30'd229266819;
array2[2588]=30'd229266819;
array2[2589]=30'd229266819;
array2[2590]=30'd231362949;
array2[2591]=30'd231362949;
array2[2592]=30'd713202349;
array2[2593]=30'd728897252;
array2[2594]=30'd718417640;
array2[2595]=30'd718417640;
array2[2596]=30'd718417640;
array2[2597]=30'd718417640;
array2[2598]=30'd718417640;
array2[2599]=30'd718417640;
array2[2600]=30'd718417640;
array2[2601]=30'd718417640;
array2[2602]=30'd672324351;
array2[2603]=30'd718417640;
array2[2604]=30'd718417640;
array2[2605]=30'd718417640;
array2[2606]=30'd728897252;
array2[2607]=30'd728897252;
array2[2608]=30'd728897252;
array2[2609]=30'd758240964;
array2[2610]=30'd728897252;
array2[2611]=30'd728897252;
array2[2612]=30'd728897252;
array2[2613]=30'd728897252;
array2[2614]=30'd728897252;
array2[2615]=30'd728897252;
array2[2616]=30'd728897252;
array2[2617]=30'd718417640;
array2[2618]=30'd718417640;
array2[2619]=30'd718417640;
array2[2620]=30'd718417640;
array2[2621]=30'd718417640;
array2[2622]=30'd672324351;
array2[2623]=30'd672324351;
array2[2624]=30'd718417640;
array2[2625]=30'd672324351;
array2[2626]=30'd672324351;
array2[2627]=30'd539218630;
array2[2628]=30'd375721588;
array2[2629]=30'd357913199;
array2[2630]=30'd606320275;
array2[2631]=30'd518272648;
array2[2632]=30'd606320275;
array2[2633]=30'd518272648;
array2[2634]=30'd672348794;
array2[2635]=30'd770812573;
array2[2636]=30'd631447172;
array2[2637]=30'd481587821;
array2[2638]=30'd481587821;
array2[2639]=30'd481587821;
array2[2640]=30'd727851632;
array2[2641]=30'd865130113;
array2[2642]=30'd858839683;
array2[2643]=30'd858839683;
array2[2644]=30'd865130113;
array2[2645]=30'd851505800;
array2[2646]=30'd565444213;
array2[2647]=30'd434416250;
array2[2648]=30'd434416250;
array2[2649]=30'd768729747;
array2[2650]=30'd851505800;
array2[2651]=30'd858839683;
array2[2652]=30'd851505800;
array2[2653]=30'd828452495;
array2[2654]=30'd819020415;
array2[2655]=30'd828452495;
array2[2656]=30'd828452495;
array2[2657]=30'd828452495;
array2[2658]=30'd851505800;
array2[2659]=30'd851505800;
array2[2660]=30'd858839683;
array2[2661]=30'd851505800;
array2[2662]=30'd851505800;
array2[2663]=30'd858839683;
array2[2664]=30'd828452495;
array2[2665]=30'd713202349;
array2[2666]=30'd461700935;
array2[2667]=30'd558174979;
array2[2668]=30'd539218630;
array2[2669]=30'd518272648;
array2[2670]=30'd677571193;
array2[2671]=30'd737318494;
array2[2672]=30'd708987491;
array2[2673]=30'd566515308;
array2[2674]=30'd319215128;
array2[2675]=30'd193577377;
array2[2676]=30'd228216193;
array2[2677]=30'd227165569;
array2[2678]=30'd231364996;
array2[2679]=30'd231362949;
array2[2680]=30'd231362949;
array2[2681]=30'd231362949;
array2[2682]=30'd230317442;
array2[2683]=30'd231362949;
array2[2684]=30'd229266819;
array2[2685]=30'd231362949;
array2[2686]=30'd229266819;
array2[2687]=30'd229266819;
array2[2688]=30'd713202349;
array2[2689]=30'd758240964;
array2[2690]=30'd718417640;
array2[2691]=30'd728897252;
array2[2692]=30'd728897252;
array2[2693]=30'd728897252;
array2[2694]=30'd728897252;
array2[2695]=30'd728897252;
array2[2696]=30'd728897252;
array2[2697]=30'd728897252;
array2[2698]=30'd728897252;
array2[2699]=30'd728897252;
array2[2700]=30'd728897252;
array2[2701]=30'd728897252;
array2[2702]=30'd728897252;
array2[2703]=30'd728897252;
array2[2704]=30'd728897252;
array2[2705]=30'd718417640;
array2[2706]=30'd728897252;
array2[2707]=30'd728897252;
array2[2708]=30'd728897252;
array2[2709]=30'd728897252;
array2[2710]=30'd728897252;
array2[2711]=30'd728897252;
array2[2712]=30'd728897252;
array2[2713]=30'd728897252;
array2[2714]=30'd728897252;
array2[2715]=30'd728897252;
array2[2716]=30'd728897252;
array2[2717]=30'd718417640;
array2[2718]=30'd728897252;
array2[2719]=30'd728897252;
array2[2720]=30'd728897252;
array2[2721]=30'd728897252;
array2[2722]=30'd728897252;
array2[2723]=30'd606320275;
array2[2724]=30'd338018898;
array2[2725]=30'd434416250;
array2[2726]=30'd331763301;
array2[2727]=30'd357913199;
array2[2728]=30'd483727963;
array2[2729]=30'd727851632;
array2[2730]=30'd828452495;
array2[2731]=30'd851505800;
array2[2732]=30'd805398138;
array2[2733]=30'd481587821;
array2[2734]=30'd481587821;
array2[2735]=30'd481587821;
array2[2736]=30'd727851632;
array2[2737]=30'd865130113;
array2[2738]=30'd858839683;
array2[2739]=30'd858839683;
array2[2740]=30'd865130113;
array2[2741]=30'd858839683;
array2[2742]=30'd764529268;
array2[2743]=30'd518272648;
array2[2744]=30'd518272648;
array2[2745]=30'd819020415;
array2[2746]=30'd851505800;
array2[2747]=30'd858839683;
array2[2748]=30'd858839683;
array2[2749]=30'd858839683;
array2[2750]=30'd865130113;
array2[2751]=30'd851505800;
array2[2752]=30'd858839683;
array2[2753]=30'd851505800;
array2[2754]=30'd851505800;
array2[2755]=30'd858839683;
array2[2756]=30'd858839683;
array2[2757]=30'd858839683;
array2[2758]=30'd865130113;
array2[2759]=30'd858839683;
array2[2760]=30'd678602388;
array2[2761]=30'd539218630;
array2[2762]=30'd537140990;
array2[2763]=30'd409311115;
array2[2764]=30'd558174979;
array2[2765]=30'd678602388;
array2[2766]=30'd737318494;
array2[2767]=30'd729975381;
array2[2768]=30'd729975381;
array2[2769]=30'd678604396;
array2[2770]=30'd506770009;
array2[2771]=30'd193577377;
array2[2772]=30'd228216193;
array2[2773]=30'd229266819;
array2[2774]=30'd231364996;
array2[2775]=30'd231364996;
array2[2776]=30'd231362949;
array2[2777]=30'd234504581;
array2[2778]=30'd229266819;
array2[2779]=30'd229266819;
array2[2780]=30'd229266819;
array2[2781]=30'd230317442;
array2[2782]=30'd231362949;
array2[2783]=30'd231362949;
array2[2784]=30'd790726247;
array2[2785]=30'd865130113;
array2[2786]=30'd799112870;
array2[2787]=30'd758240964;
array2[2788]=30'd728897252;
array2[2789]=30'd728897252;
array2[2790]=30'd728897252;
array2[2791]=30'd728897252;
array2[2792]=30'd728897252;
array2[2793]=30'd728897252;
array2[2794]=30'd728897252;
array2[2795]=30'd728897252;
array2[2796]=30'd728897252;
array2[2797]=30'd758240964;
array2[2798]=30'd865130113;
array2[2799]=30'd851505800;
array2[2800]=30'd865130113;
array2[2801]=30'd858839683;
array2[2802]=30'd865130113;
array2[2803]=30'd858839683;
array2[2804]=30'd858839683;
array2[2805]=30'd865130113;
array2[2806]=30'd858839683;
array2[2807]=30'd865130113;
array2[2808]=30'd865130113;
array2[2809]=30'd851505800;
array2[2810]=30'd758240964;
array2[2811]=30'd728897252;
array2[2812]=30'd728897252;
array2[2813]=30'd728897252;
array2[2814]=30'd718417640;
array2[2815]=30'd728897252;
array2[2816]=30'd718417640;
array2[2817]=30'd728897252;
array2[2818]=30'd728897252;
array2[2819]=30'd606320275;
array2[2820]=30'd299264555;
array2[2821]=30'd347490866;
array2[2822]=30'd265736724;
array2[2823]=30'd434416250;
array2[2824]=30'd713179821;
array2[2825]=30'd828452495;
array2[2826]=30'd851505800;
array2[2827]=30'd858839683;
array2[2828]=30'd851505800;
array2[2829]=30'd678602388;
array2[2830]=30'd481587821;
array2[2831]=30'd481587821;
array2[2832]=30'd727851632;
array2[2833]=30'd865130113;
array2[2834]=30'd858839683;
array2[2835]=30'd858839683;
array2[2836]=30'd865130113;
array2[2837]=30'd858839683;
array2[2838]=30'd851505800;
array2[2839]=30'd768729747;
array2[2840]=30'd764529268;
array2[2841]=30'd851505800;
array2[2842]=30'd858839683;
array2[2843]=30'd865130113;
array2[2844]=30'd858839683;
array2[2845]=30'd858839683;
array2[2846]=30'd865130113;
array2[2847]=30'd865130113;
array2[2848]=30'd858839683;
array2[2849]=30'd858839683;
array2[2850]=30'd865130113;
array2[2851]=30'd858839683;
array2[2852]=30'd865130113;
array2[2853]=30'd858839683;
array2[2854]=30'd865130113;
array2[2855]=30'd851505800;
array2[2856]=30'd601041592;
array2[2857]=30'd451191548;
array2[2858]=30'd451191548;
array2[2859]=30'd390446940;
array2[2860]=30'd461700935;
array2[2861]=30'd646169309;
array2[2862]=30'd737318494;
array2[2863]=30'd737318494;
array2[2864]=30'd708987491;
array2[2865]=30'd566515308;
array2[2866]=30'd383147560;
array2[2867]=30'd207191473;
array2[2868]=30'd231359873;
array2[2869]=30'd229266819;
array2[2870]=30'd231362949;
array2[2871]=30'd229266819;
array2[2872]=30'd231362949;
array2[2873]=30'd229266819;
array2[2874]=30'd231362949;
array2[2875]=30'd231359873;
array2[2876]=30'd231362949;
array2[2877]=30'd231364996;
array2[2878]=30'd231364996;
array2[2879]=30'd231362949;
array2[2880]=30'd823228019;
array2[2881]=30'd906004072;
array2[2882]=30'd906004072;
array2[2883]=30'd865130113;
array2[2884]=30'd865130113;
array2[2885]=30'd865130113;
array2[2886]=30'd865130113;
array2[2887]=30'd865130113;
array2[2888]=30'd858839683;
array2[2889]=30'd865130113;
array2[2890]=30'd865130113;
array2[2891]=30'd865130113;
array2[2892]=30'd865130113;
array2[2893]=30'd865130113;
array2[2894]=30'd906004072;
array2[2895]=30'd906004072;
array2[2896]=30'd906004072;
array2[2897]=30'd906004072;
array2[2898]=30'd906004072;
array2[2899]=30'd906004072;
array2[2900]=30'd906004072;
array2[2901]=30'd906004072;
array2[2902]=30'd906004072;
array2[2903]=30'd906004072;
array2[2904]=30'd906004072;
array2[2905]=30'd906004072;
array2[2906]=30'd865130113;
array2[2907]=30'd865130113;
array2[2908]=30'd865130113;
array2[2909]=30'd865130113;
array2[2910]=30'd865130113;
array2[2911]=30'd865130113;
array2[2912]=30'd865130113;
array2[2913]=30'd865130113;
array2[2914]=30'd865130113;
array2[2915]=30'd819020415;
array2[2916]=30'd790726247;
array2[2917]=30'd790726247;
array2[2918]=30'd678604396;
array2[2919]=30'd407216718;
array2[2920]=30'd828452495;
array2[2921]=30'd851505800;
array2[2922]=30'd858839683;
array2[2923]=30'd851505800;
array2[2924]=30'd858839683;
array2[2925]=30'd828452495;
array2[2926]=30'd678602388;
array2[2927]=30'd481587821;
array2[2928]=30'd727851632;
array2[2929]=30'd858839683;
array2[2930]=30'd865130113;
array2[2931]=30'd858839683;
array2[2932]=30'd851505800;
array2[2933]=30'd865130113;
array2[2934]=30'd865130113;
array2[2935]=30'd858839683;
array2[2936]=30'd865130113;
array2[2937]=30'd865130113;
array2[2938]=30'd858839683;
array2[2939]=30'd865130113;
array2[2940]=30'd865130113;
array2[2941]=30'd858839683;
array2[2942]=30'd858839683;
array2[2943]=30'd858839683;
array2[2944]=30'd865130113;
array2[2945]=30'd858839683;
array2[2946]=30'd858839683;
array2[2947]=30'd865130113;
array2[2948]=30'd858839683;
array2[2949]=30'd865130113;
array2[2950]=30'd858839683;
array2[2951]=30'd858839683;
array2[2952]=30'd770812573;
array2[2953]=30'd601041592;
array2[2954]=30'd395649781;
array2[2955]=30'd395649781;
array2[2956]=30'd601041592;
array2[2957]=30'd727851632;
array2[2958]=30'd727851632;
array2[2959]=30'd729975381;
array2[2960]=30'd708987491;
array2[2961]=30'd538207812;
array2[2962]=30'd195647926;
array2[2963]=30'd210373000;
array2[2964]=30'd231364996;
array2[2965]=30'd229266819;
array2[2966]=30'd229266819;
array2[2967]=30'd231364996;
array2[2968]=30'd229266819;
array2[2969]=30'd231362949;
array2[2970]=30'd231362949;
array2[2971]=30'd231362949;
array2[2972]=30'd231362949;
array2[2973]=30'd229266819;
array2[2974]=30'd231364996;
array2[2975]=30'd231362949;
array2[2976]=30'd823228019;
array2[2977]=30'd906004072;
array2[2978]=30'd906004072;
array2[2979]=30'd906004072;
array2[2980]=30'd906004072;
array2[2981]=30'd906004072;
array2[2982]=30'd906004072;
array2[2983]=30'd906004072;
array2[2984]=30'd906004072;
array2[2985]=30'd906004072;
array2[2986]=30'd906004072;
array2[2987]=30'd906004072;
array2[2988]=30'd906004072;
array2[2989]=30'd906004072;
array2[2990]=30'd906004072;
array2[2991]=30'd906004072;
array2[2992]=30'd906004072;
array2[2993]=30'd906004072;
array2[2994]=30'd906004072;
array2[2995]=30'd906004072;
array2[2996]=30'd906004072;
array2[2997]=30'd906004072;
array2[2998]=30'd906004072;
array2[2999]=30'd906004072;
array2[3000]=30'd906004072;
array2[3001]=30'd906004072;
array2[3002]=30'd906004072;
array2[3003]=30'd906004072;
array2[3004]=30'd906004072;
array2[3005]=30'd906004072;
array2[3006]=30'd906004072;
array2[3007]=30'd906004072;
array2[3008]=30'd906004072;
array2[3009]=30'd906004072;
array2[3010]=30'd906004072;
array2[3011]=30'd906004072;
array2[3012]=30'd906004072;
array2[3013]=30'd906004072;
array2[3014]=30'd678604396;
array2[3015]=30'd483727963;
array2[3016]=30'd865130113;
array2[3017]=30'd865130113;
array2[3018]=30'd858839683;
array2[3019]=30'd858839683;
array2[3020]=30'd865130113;
array2[3021]=30'd858839683;
array2[3022]=30'd828452495;
array2[3023]=30'd677571193;
array2[3024]=30'd762499681;
array2[3025]=30'd858839683;
array2[3026]=30'd858839683;
array2[3027]=30'd858839683;
array2[3028]=30'd865130113;
array2[3029]=30'd858839683;
array2[3030]=30'd858839683;
array2[3031]=30'd865130113;
array2[3032]=30'd865130113;
array2[3033]=30'd858839683;
array2[3034]=30'd858839683;
array2[3035]=30'd865130113;
array2[3036]=30'd858839683;
array2[3037]=30'd858839683;
array2[3038]=30'd858839683;
array2[3039]=30'd865130113;
array2[3040]=30'd858839683;
array2[3041]=30'd858839683;
array2[3042]=30'd865130113;
array2[3043]=30'd865130113;
array2[3044]=30'd828452495;
array2[3045]=30'd819020415;
array2[3046]=30'd828452495;
array2[3047]=30'd851505800;
array2[3048]=30'd828452495;
array2[3049]=30'd770812573;
array2[3050]=30'd451191548;
array2[3051]=30'd537140990;
array2[3052]=30'd770812573;
array2[3053]=30'd764529268;
array2[3054]=30'd727851632;
array2[3055]=30'd678604396;
array2[3056]=30'd645112409;
array2[3057]=30'd401997362;
array2[3058]=30'd207191473;
array2[3059]=30'd231359873;
array2[3060]=30'd231364996;
array2[3061]=30'd231362949;
array2[3062]=30'd229266819;
array2[3063]=30'd230317442;
array2[3064]=30'd231364996;
array2[3065]=30'd228216193;
array2[3066]=30'd231362949;
array2[3067]=30'd234504581;
array2[3068]=30'd229266819;
array2[3069]=30'd229266819;
array2[3070]=30'd229266819;
array2[3071]=30'd229266819;
array2[3072]=30'd736232864;
array2[3073]=30'd690121052;
array2[3074]=30'd783393281;
array2[3075]=30'd906004072;
array2[3076]=30'd906004072;
array2[3077]=30'd906004072;
array2[3078]=30'd906004072;
array2[3079]=30'd906004072;
array2[3080]=30'd906004072;
array2[3081]=30'd906004072;
array2[3082]=30'd906004072;
array2[3083]=30'd906004072;
array2[3084]=30'd906004072;
array2[3085]=30'd832648722;
array2[3086]=30'd690121052;
array2[3087]=30'd690121052;
array2[3088]=30'd690121052;
array2[3089]=30'd690121052;
array2[3090]=30'd690121052;
array2[3091]=30'd690121052;
array2[3092]=30'd690121052;
array2[3093]=30'd690121052;
array2[3094]=30'd690121052;
array2[3095]=30'd690121052;
array2[3096]=30'd690121052;
array2[3097]=30'd736232864;
array2[3098]=30'd906004072;
array2[3099]=30'd906004072;
array2[3100]=30'd906004072;
array2[3101]=30'd906004072;
array2[3102]=30'd906004072;
array2[3103]=30'd906004072;
array2[3104]=30'd906004072;
array2[3105]=30'd906004072;
array2[3106]=30'd906004072;
array2[3107]=30'd906004072;
array2[3108]=30'd823228019;
array2[3109]=30'd736232864;
array2[3110]=30'd352736774;
array2[3111]=30'd764529268;
array2[3112]=30'd851505800;
array2[3113]=30'd858839683;
array2[3114]=30'd858839683;
array2[3115]=30'd858839683;
array2[3116]=30'd858839683;
array2[3117]=30'd865130113;
array2[3118]=30'd858839683;
array2[3119]=30'd858839683;
array2[3120]=30'd858839683;
array2[3121]=30'd858839683;
array2[3122]=30'd858839683;
array2[3123]=30'd858839683;
array2[3124]=30'd858839683;
array2[3125]=30'd858839683;
array2[3126]=30'd858839683;
array2[3127]=30'd858839683;
array2[3128]=30'd858839683;
array2[3129]=30'd858839683;
array2[3130]=30'd858839683;
array2[3131]=30'd858839683;
array2[3132]=30'd858839683;
array2[3133]=30'd865130113;
array2[3134]=30'd858839683;
array2[3135]=30'd858839683;
array2[3136]=30'd858839683;
array2[3137]=30'd865130113;
array2[3138]=30'd865130113;
array2[3139]=30'd858839683;
array2[3140]=30'd711090860;
array2[3141]=30'd606320275;
array2[3142]=30'd678602388;
array2[3143]=30'd713179821;
array2[3144]=30'd732038833;
array2[3145]=30'd770812573;
array2[3146]=30'd678602388;
array2[3147]=30'd678602388;
array2[3148]=30'd770812573;
array2[3149]=30'd678602388;
array2[3150]=30'd631447172;
array2[3151]=30'd631447172;
array2[3152]=30'd444954173;
array2[3153]=30'd195647926;
array2[3154]=30'd227159434;
array2[3155]=30'd231362949;
array2[3156]=30'd231362949;
array2[3157]=30'd230317442;
array2[3158]=30'd229266819;
array2[3159]=30'd231362949;
array2[3160]=30'd228216193;
array2[3161]=30'd227165569;
array2[3162]=30'd231362949;
array2[3163]=30'd231359873;
array2[3164]=30'd229266819;
array2[3165]=30'd230317442;
array2[3166]=30'd229266819;
array2[3167]=30'd231362949;
array2[3168]=30'd582318295;
array2[3169]=30'd611520752;
array2[3170]=30'd637725975;
array2[3171]=30'd690121052;
array2[3172]=30'd690121052;
array2[3173]=30'd690121052;
array2[3174]=30'd690121052;
array2[3175]=30'd690121052;
array2[3176]=30'd690121052;
array2[3177]=30'd736232864;
array2[3178]=30'd690121052;
array2[3179]=30'd736232864;
array2[3180]=30'd736232864;
array2[3181]=30'd690121052;
array2[3182]=30'd611520752;
array2[3183]=30'd611520752;
array2[3184]=30'd611520752;
array2[3185]=30'd611520752;
array2[3186]=30'd611520752;
array2[3187]=30'd611520752;
array2[3188]=30'd611520752;
array2[3189]=30'd606284005;
array2[3190]=30'd611520752;
array2[3191]=30'd611520752;
array2[3192]=30'd606284005;
array2[3193]=30'd615715061;
array2[3194]=30'd690121052;
array2[3195]=30'd736232864;
array2[3196]=30'd736232864;
array2[3197]=30'd736232864;
array2[3198]=30'd690121052;
array2[3199]=30'd736232864;
array2[3200]=30'd736232864;
array2[3201]=30'd690121052;
array2[3202]=30'd690121052;
array2[3203]=30'd736232864;
array2[3204]=30'd690121052;
array2[3205]=30'd619916568;
array2[3206]=30'd281508345;
array2[3207]=30'd819020415;
array2[3208]=30'd828452495;
array2[3209]=30'd851505800;
array2[3210]=30'd865130113;
array2[3211]=30'd858839683;
array2[3212]=30'd858839683;
array2[3213]=30'd865130113;
array2[3214]=30'd858839683;
array2[3215]=30'd858839683;
array2[3216]=30'd865130113;
array2[3217]=30'd865130113;
array2[3218]=30'd858839683;
array2[3219]=30'd858839683;
array2[3220]=30'd865130113;
array2[3221]=30'd858839683;
array2[3222]=30'd858839683;
array2[3223]=30'd865130113;
array2[3224]=30'd858839683;
array2[3225]=30'd858839683;
array2[3226]=30'd858839683;
array2[3227]=30'd865130113;
array2[3228]=30'd865130113;
array2[3229]=30'd858839683;
array2[3230]=30'd858839683;
array2[3231]=30'd858839683;
array2[3232]=30'd865130113;
array2[3233]=30'd858839683;
array2[3234]=30'd858839683;
array2[3235]=30'd865130113;
array2[3236]=30'd851505800;
array2[3237]=30'd770812573;
array2[3238]=30'd672348794;
array2[3239]=30'd672348794;
array2[3240]=30'd606320275;
array2[3241]=30'd678602388;
array2[3242]=30'd601041592;
array2[3243]=30'd711090860;
array2[3244]=30'd770812573;
array2[3245]=30'd678602388;
array2[3246]=30'd566515308;
array2[3247]=30'd407216718;
array2[3248]=30'd195647926;
array2[3249]=30'd230307208;
array2[3250]=30'd234504581;
array2[3251]=30'd231362949;
array2[3252]=30'd230317442;
array2[3253]=30'd228212100;
array2[3254]=30'd228216193;
array2[3255]=30'd229266819;
array2[3256]=30'd230317442;
array2[3257]=30'd231364996;
array2[3258]=30'd231362949;
array2[3259]=30'd234504581;
array2[3260]=30'd229266819;
array2[3261]=30'd231362949;
array2[3262]=30'd229266819;
array2[3263]=30'd230317442;
array2[3264]=30'd582318295;
array2[3265]=30'd611520752;
array2[3266]=30'd606284005;
array2[3267]=30'd606284005;
array2[3268]=30'd611520752;
array2[3269]=30'd606284005;
array2[3270]=30'd606284005;
array2[3271]=30'd606284005;
array2[3272]=30'd611520752;
array2[3273]=30'd606284005;
array2[3274]=30'd606284005;
array2[3275]=30'd606284005;
array2[3276]=30'd611520752;
array2[3277]=30'd606284005;
array2[3278]=30'd611520752;
array2[3279]=30'd606284005;
array2[3280]=30'd611520752;
array2[3281]=30'd606284005;
array2[3282]=30'd611520752;
array2[3283]=30'd611520752;
array2[3284]=30'd606284005;
array2[3285]=30'd611520752;
array2[3286]=30'd611520752;
array2[3287]=30'd611520752;
array2[3288]=30'd611520752;
array2[3289]=30'd611520752;
array2[3290]=30'd606284005;
array2[3291]=30'd611520752;
array2[3292]=30'd611520752;
array2[3293]=30'd606284005;
array2[3294]=30'd611520752;
array2[3295]=30'd606284005;
array2[3296]=30'd606284005;
array2[3297]=30'd606284005;
array2[3298]=30'd611520752;
array2[3299]=30'd611520752;
array2[3300]=30'd611520752;
array2[3301]=30'd521469272;
array2[3302]=30'd538207812;
array2[3303]=30'd851505800;
array2[3304]=30'd858839683;
array2[3305]=30'd858839683;
array2[3306]=30'd858839683;
array2[3307]=30'd865130113;
array2[3308]=30'd865130113;
array2[3309]=30'd858839683;
array2[3310]=30'd865130113;
array2[3311]=30'd865130113;
array2[3312]=30'd858839683;
array2[3313]=30'd858839683;
array2[3314]=30'd858839683;
array2[3315]=30'd865130113;
array2[3316]=30'd865130113;
array2[3317]=30'd858839683;
array2[3318]=30'd858839683;
array2[3319]=30'd865130113;
array2[3320]=30'd858839683;
array2[3321]=30'd858839683;
array2[3322]=30'd858839683;
array2[3323]=30'd865130113;
array2[3324]=30'd865130113;
array2[3325]=30'd858839683;
array2[3326]=30'd858839683;
array2[3327]=30'd865130113;
array2[3328]=30'd858839683;
array2[3329]=30'd865130113;
array2[3330]=30'd865130113;
array2[3331]=30'd858839683;
array2[3332]=30'd828452495;
array2[3333]=30'd799112870;
array2[3334]=30'd758240964;
array2[3335]=30'd799112870;
array2[3336]=30'd711090860;
array2[3337]=30'd678602388;
array2[3338]=30'd560184961;
array2[3339]=30'd604201637;
array2[3340]=30'd631447172;
array2[3341]=30'd560184961;
array2[3342]=30'd434416250;
array2[3343]=30'd338018898;
array2[3344]=30'd195647926;
array2[3345]=30'd212454818;
array2[3346]=30'd227165569;
array2[3347]=30'd229266819;
array2[3348]=30'd230317442;
array2[3349]=30'd230317442;
array2[3350]=30'd228216193;
array2[3351]=30'd231362949;
array2[3352]=30'd231362949;
array2[3353]=30'd229266819;
array2[3354]=30'd229266819;
array2[3355]=30'd229266819;
array2[3356]=30'd229266819;
array2[3357]=30'd231362949;
array2[3358]=30'd231362949;
array2[3359]=30'd234504581;
array2[3360]=30'd559433927;
array2[3361]=30'd585627858;
array2[3362]=30'd586531028;
array2[3363]=30'd606284005;
array2[3364]=30'd606284005;
array2[3365]=30'd606284005;
array2[3366]=30'd611520752;
array2[3367]=30'd606284005;
array2[3368]=30'd611520752;
array2[3369]=30'd606284005;
array2[3370]=30'd611520752;
array2[3371]=30'd606284005;
array2[3372]=30'd606284005;
array2[3373]=30'd595854564;
array2[3374]=30'd585627858;
array2[3375]=30'd585627858;
array2[3376]=30'd585627858;
array2[3377]=30'd585627858;
array2[3378]=30'd585627858;
array2[3379]=30'd585627858;
array2[3380]=30'd585627858;
array2[3381]=30'd585627858;
array2[3382]=30'd585627858;
array2[3383]=30'd585627858;
array2[3384]=30'd585627858;
array2[3385]=30'd585627858;
array2[3386]=30'd606284005;
array2[3387]=30'd606284005;
array2[3388]=30'd606284005;
array2[3389]=30'd606284005;
array2[3390]=30'd606284005;
array2[3391]=30'd606284005;
array2[3392]=30'd606284005;
array2[3393]=30'd606284005;
array2[3394]=30'd611520752;
array2[3395]=30'd606284005;
array2[3396]=30'd606284005;
array2[3397]=30'd281508345;
array2[3398]=30'd678602388;
array2[3399]=30'd851505800;
array2[3400]=30'd865130113;
array2[3401]=30'd858839683;
array2[3402]=30'd851505800;
array2[3403]=30'd865130113;
array2[3404]=30'd858839683;
array2[3405]=30'd858839683;
array2[3406]=30'd858839683;
array2[3407]=30'd865130113;
array2[3408]=30'd865130113;
array2[3409]=30'd865130113;
array2[3410]=30'd858839683;
array2[3411]=30'd858839683;
array2[3412]=30'd865130113;
array2[3413]=30'd858839683;
array2[3414]=30'd865130113;
array2[3415]=30'd858839683;
array2[3416]=30'd865130113;
array2[3417]=30'd858839683;
array2[3418]=30'd858839683;
array2[3419]=30'd865130113;
array2[3420]=30'd858839683;
array2[3421]=30'd858839683;
array2[3422]=30'd865130113;
array2[3423]=30'd865130113;
array2[3424]=30'd858839683;
array2[3425]=30'd851505800;
array2[3426]=30'd858839683;
array2[3427]=30'd851505800;
array2[3428]=30'd770812573;
array2[3429]=30'd770812573;
array2[3430]=30'd770812573;
array2[3431]=30'd770812573;
array2[3432]=30'd799112870;
array2[3433]=30'd828452495;
array2[3434]=30'd768729747;
array2[3435]=30'd678602388;
array2[3436]=30'd566515308;
array2[3437]=30'd566515308;
array2[3438]=30'd606320275;
array2[3439]=30'd485780117;
array2[3440]=30'd449120871;
array2[3441]=30'd319215128;
array2[3442]=30'd212454818;
array2[3443]=30'd228216193;
array2[3444]=30'd228216193;
array2[3445]=30'd231364996;
array2[3446]=30'd231364996;
array2[3447]=30'd231362949;
array2[3448]=30'd231362949;
array2[3449]=30'd231359873;
array2[3450]=30'd229266819;
array2[3451]=30'd229266819;
array2[3452]=30'd229266819;
array2[3453]=30'd229266819;
array2[3454]=30'd231362949;
array2[3455]=30'd231362949;
array2[3456]=30'd530274492;
array2[3457]=30'd524037312;
array2[3458]=30'd530274492;
array2[3459]=30'd561572038;
array2[3460]=30'd561572038;
array2[3461]=30'd561572038;
array2[3462]=30'd561572038;
array2[3463]=30'd561572038;
array2[3464]=30'd561572038;
array2[3465]=30'd561572038;
array2[3466]=30'd561572038;
array2[3467]=30'd561572038;
array2[3468]=30'd561572038;
array2[3469]=30'd543866052;
array2[3470]=30'd524037312;
array2[3471]=30'd518815920;
array2[3472]=30'd518815920;
array2[3473]=30'd518815920;
array2[3474]=30'd518815920;
array2[3475]=30'd518815920;
array2[3476]=30'd518815920;
array2[3477]=30'd518815920;
array2[3478]=30'd518815920;
array2[3479]=30'd518815920;
array2[3480]=30'd518815920;
array2[3481]=30'd514590904;
array2[3482]=30'd561572038;
array2[3483]=30'd561572038;
array2[3484]=30'd561572038;
array2[3485]=30'd561572038;
array2[3486]=30'd561572038;
array2[3487]=30'd561572038;
array2[3488]=30'd561572038;
array2[3489]=30'd561572038;
array2[3490]=30'd561572038;
array2[3491]=30'd561572038;
array2[3492]=30'd543866052;
array2[3493]=30'd304706973;
array2[3494]=30'd727851632;
array2[3495]=30'd828452495;
array2[3496]=30'd865130113;
array2[3497]=30'd858839683;
array2[3498]=30'd851505800;
array2[3499]=30'd858839683;
array2[3500]=30'd865130113;
array2[3501]=30'd858839683;
array2[3502]=30'd858839683;
array2[3503]=30'd865130113;
array2[3504]=30'd865130113;
array2[3505]=30'd858839683;
array2[3506]=30'd851505800;
array2[3507]=30'd851505800;
array2[3508]=30'd851505800;
array2[3509]=30'd851505800;
array2[3510]=30'd851505800;
array2[3511]=30'd851505800;
array2[3512]=30'd858839683;
array2[3513]=30'd858839683;
array2[3514]=30'd865130113;
array2[3515]=30'd858839683;
array2[3516]=30'd858839683;
array2[3517]=30'd851505800;
array2[3518]=30'd851505800;
array2[3519]=30'd799112870;
array2[3520]=30'd770812573;
array2[3521]=30'd768729747;
array2[3522]=30'd770812573;
array2[3523]=30'd770812573;
array2[3524]=30'd732038833;
array2[3525]=30'd770812573;
array2[3526]=30'd770812573;
array2[3527]=30'd770812573;
array2[3528]=30'd799112870;
array2[3529]=30'd828452495;
array2[3530]=30'd851505800;
array2[3531]=30'd851505800;
array2[3532]=30'd770816666;
array2[3533]=30'd631447172;
array2[3534]=30'd566515308;
array2[3535]=30'd434416250;
array2[3536]=30'd407216718;
array2[3537]=30'd260631016;
array2[3538]=30'd232392085;
array2[3539]=30'd227165569;
array2[3540]=30'd231362949;
array2[3541]=30'd229266819;
array2[3542]=30'd231364996;
array2[3543]=30'd231359873;
array2[3544]=30'd229266819;
array2[3545]=30'd229266819;
array2[3546]=30'd231359873;
array2[3547]=30'd231362949;
array2[3548]=30'd231362949;
array2[3549]=30'd231364996;
array2[3550]=30'd231362949;
array2[3551]=30'd231362949;
array2[3552]=30'd518785242;
array2[3553]=30'd518815920;
array2[3554]=30'd521966763;
array2[3555]=30'd521966763;
array2[3556]=30'd518815920;
array2[3557]=30'd521966763;
array2[3558]=30'd518815920;
array2[3559]=30'd518815920;
array2[3560]=30'd518815920;
array2[3561]=30'd518815920;
array2[3562]=30'd518815920;
array2[3563]=30'd518815920;
array2[3564]=30'd521966763;
array2[3565]=30'd521966763;
array2[3566]=30'd521966763;
array2[3567]=30'd521966763;
array2[3568]=30'd521966763;
array2[3569]=30'd521966763;
array2[3570]=30'd521966763;
array2[3571]=30'd521966763;
array2[3572]=30'd521966763;
array2[3573]=30'd521966763;
array2[3574]=30'd518815920;
array2[3575]=30'd521966763;
array2[3576]=30'd521966763;
array2[3577]=30'd521966763;
array2[3578]=30'd521966763;
array2[3579]=30'd521966763;
array2[3580]=30'd518815920;
array2[3581]=30'd518815920;
array2[3582]=30'd518815920;
array2[3583]=30'd521966763;
array2[3584]=30'd521966763;
array2[3585]=30'd521966763;
array2[3586]=30'd521966763;
array2[3587]=30'd518815920;
array2[3588]=30'd521966763;
array2[3589]=30'd338288022;
array2[3590]=30'd678602388;
array2[3591]=30'd851505800;
array2[3592]=30'd851505800;
array2[3593]=30'd858839683;
array2[3594]=30'd858839683;
array2[3595]=30'd858839683;
array2[3596]=30'd858839683;
array2[3597]=30'd851505800;
array2[3598]=30'd819020415;
array2[3599]=30'd828452495;
array2[3600]=30'd851505800;
array2[3601]=30'd851505800;
array2[3602]=30'd851505800;
array2[3603]=30'd851505800;
array2[3604]=30'd851505800;
array2[3605]=30'd851505800;
array2[3606]=30'd828452495;
array2[3607]=30'd828452495;
array2[3608]=30'd828452495;
array2[3609]=30'd828452495;
array2[3610]=30'd851505800;
array2[3611]=30'd799112870;
array2[3612]=30'd799112870;
array2[3613]=30'd799112870;
array2[3614]=30'd770812573;
array2[3615]=30'd711090860;
array2[3616]=30'd631447172;
array2[3617]=30'd506770009;
array2[3618]=30'd631447172;
array2[3619]=30'd678602388;
array2[3620]=30'd713179821;
array2[3621]=30'd713202349;
array2[3622]=30'd713202349;
array2[3623]=30'd732038833;
array2[3624]=30'd799112870;
array2[3625]=30'd851505800;
array2[3626]=30'd851505800;
array2[3627]=30'd858839683;
array2[3628]=30'd851505800;
array2[3629]=30'd770812573;
array2[3630]=30'd631447172;
array2[3631]=30'd401997362;
array2[3632]=30'd190356956;
array2[3633]=30'd220861839;
array2[3634]=30'd229266819;
array2[3635]=30'd231362949;
array2[3636]=30'd230317442;
array2[3637]=30'd231364996;
array2[3638]=30'd231362949;
array2[3639]=30'd231362949;
array2[3640]=30'd231359873;
array2[3641]=30'd229266819;
array2[3642]=30'd229266819;
array2[3643]=30'd229266819;
array2[3644]=30'd229266819;
array2[3645]=30'd231362949;
array2[3646]=30'd231362949;
array2[3647]=30'd234504581;
array2[3648]=30'd520893723;
array2[3649]=30'd510427417;
array2[3650]=30'd515671261;
array2[3651]=30'd518815920;
array2[3652]=30'd521966763;
array2[3653]=30'd518815920;
array2[3654]=30'd521966763;
array2[3655]=30'd521966763;
array2[3656]=30'd521966763;
array2[3657]=30'd521966763;
array2[3658]=30'd521966763;
array2[3659]=30'd521966763;
array2[3660]=30'd521966763;
array2[3661]=30'd518815920;
array2[3662]=30'd510427417;
array2[3663]=30'd510427417;
array2[3664]=30'd510427417;
array2[3665]=30'd510427417;
array2[3666]=30'd510427417;
array2[3667]=30'd510427417;
array2[3668]=30'd510427417;
array2[3669]=30'd510427417;
array2[3670]=30'd510427417;
array2[3671]=30'd510427417;
array2[3672]=30'd510427417;
array2[3673]=30'd515671261;
array2[3674]=30'd518815920;
array2[3675]=30'd521966763;
array2[3676]=30'd518815920;
array2[3677]=30'd521966763;
array2[3678]=30'd521966763;
array2[3679]=30'd521966763;
array2[3680]=30'd521966763;
array2[3681]=30'd521966763;
array2[3682]=30'd518815920;
array2[3683]=30'd518815920;
array2[3684]=30'd518815920;
array2[3685]=30'd338288022;
array2[3686]=30'd711090860;
array2[3687]=30'd828452495;
array2[3688]=30'd851505800;
array2[3689]=30'd858839683;
array2[3690]=30'd858839683;
array2[3691]=30'd851505800;
array2[3692]=30'd828452495;
array2[3693]=30'd819020415;
array2[3694]=30'd768729747;
array2[3695]=30'd805398138;
array2[3696]=30'd819020415;
array2[3697]=30'd805398138;
array2[3698]=30'd805398138;
array2[3699]=30'd770816666;
array2[3700]=30'd805398138;
array2[3701]=30'd770812573;
array2[3702]=30'd799112870;
array2[3703]=30'd758240964;
array2[3704]=30'd732038833;
array2[3705]=30'd732038833;
array2[3706]=30'd758240964;
array2[3707]=30'd770812573;
array2[3708]=30'd732038833;
array2[3709]=30'd678602388;
array2[3710]=30'd631447172;
array2[3711]=30'd481587821;
array2[3712]=30'd319215128;
array2[3713]=30'd281508345;
array2[3714]=30'd281508345;
array2[3715]=30'd319215128;
array2[3716]=30'd560184961;
array2[3717]=30'd631447172;
array2[3718]=30'd601041592;
array2[3719]=30'd713202349;
array2[3720]=30'd770812573;
array2[3721]=30'd770812573;
array2[3722]=30'd799112870;
array2[3723]=30'd828452495;
array2[3724]=30'd828452495;
array2[3725]=30'd770816666;
array2[3726]=30'd565444213;
array2[3727]=30'd190356956;
array2[3728]=30'd227159434;
array2[3729]=30'd231362949;
array2[3730]=30'd231364996;
array2[3731]=30'd272255371;
array2[3732]=30'd553231776;
array2[3733]=30'd377085336;
array2[3734]=30'd227159434;
array2[3735]=30'd228216193;
array2[3736]=30'd231362949;
array2[3737]=30'd229266819;
array2[3738]=30'd231359873;
array2[3739]=30'd229266819;
array2[3740]=30'd231362949;
array2[3741]=30'd231359873;
array2[3742]=30'd231362949;
array2[3743]=30'd231362949;
array2[3744]=30'd457992679;
array2[3745]=30'd482138634;
array2[3746]=30'd477946350;
array2[3747]=30'd482131304;
array2[3748]=30'd482131304;
array2[3749]=30'd482131304;
array2[3750]=30'd482131304;
array2[3751]=30'd482131304;
array2[3752]=30'd482131304;
array2[3753]=30'd482131304;
array2[3754]=30'd482131304;
array2[3755]=30'd482131304;
array2[3756]=30'd482131304;
array2[3757]=30'd475838865;
array2[3758]=30'd477946350;
array2[3759]=30'd482138634;
array2[3760]=30'd482138634;
array2[3761]=30'd482138634;
array2[3762]=30'd482138634;
array2[3763]=30'd482138634;
array2[3764]=30'd482138634;
array2[3765]=30'd482138634;
array2[3766]=30'd480046615;
array2[3767]=30'd480046615;
array2[3768]=30'd480046615;
array2[3769]=30'd477946350;
array2[3770]=30'd475838865;
array2[3771]=30'd482131304;
array2[3772]=30'd482131304;
array2[3773]=30'd482131304;
array2[3774]=30'd482131304;
array2[3775]=30'd482131304;
array2[3776]=30'd482131304;
array2[3777]=30'd482131304;
array2[3778]=30'd482131304;
array2[3779]=30'd482131304;
array2[3780]=30'd462205301;
array2[3781]=30'd280568333;
array2[3782]=30'd711090860;
array2[3783]=30'd764529268;
array2[3784]=30'd770812573;
array2[3785]=30'd805398138;
array2[3786]=30'd805398138;
array2[3787]=30'd805398138;
array2[3788]=30'd805398138;
array2[3789]=30'd764529268;
array2[3790]=30'd737318494;
array2[3791]=30'd749877860;
array2[3792]=30'd708987491;
array2[3793]=30'd708987491;
array2[3794]=30'd672348794;
array2[3795]=30'd631447172;
array2[3796]=30'd631447172;
array2[3797]=30'd672348794;
array2[3798]=30'd711090860;
array2[3799]=30'd713179821;
array2[3800]=30'd732038833;
array2[3801]=30'd678602388;
array2[3802]=30'd606320275;
array2[3803]=30'd606320275;
array2[3804]=30'd560184961;
array2[3805]=30'd352736774;
array2[3806]=30'd281508345;
array2[3807]=30'd339244483;
array2[3808]=30'd356016571;
array2[3809]=30'd339244483;
array2[3810]=30'd339244483;
array2[3811]=30'd356016571;
array2[3812]=30'd339244483;
array2[3813]=30'd281508345;
array2[3814]=30'd401997362;
array2[3815]=30'd560184961;
array2[3816]=30'd606320275;
array2[3817]=30'd631447172;
array2[3818]=30'd631447172;
array2[3819]=30'd631447172;
array2[3820]=30'd606320275;
array2[3821]=30'd481587821;
array2[3822]=30'd347490866;
array2[3823]=30'd179916222;
array2[3824]=30'd230307208;
array2[3825]=30'd532258209;
array2[3826]=30'd377085336;
array2[3827]=30'd272255371;
array2[3828]=30'd532258209;
array2[3829]=30'd338288022;
array2[3830]=30'd338288022;
array2[3831]=30'd532258209;
array2[3832]=30'd262793620;
array2[3833]=30'd227165569;
array2[3834]=30'd231359873;
array2[3835]=30'd229266819;
array2[3836]=30'd230317442;
array2[3837]=30'd229266819;
array2[3838]=30'd234504581;
array2[3839]=30'd231362949;
array2[3840]=30'd457992679;
array2[3841]=30'd480046615;
array2[3842]=30'd480046615;
array2[3843]=30'd480046615;
array2[3844]=30'd475850257;
array2[3845]=30'd480046615;
array2[3846]=30'd480046615;
array2[3847]=30'd480046615;
array2[3848]=30'd480046615;
array2[3849]=30'd480046615;
array2[3850]=30'd480046615;
array2[3851]=30'd475850257;
array2[3852]=30'd475850257;
array2[3853]=30'd480046615;
array2[3854]=30'd480046615;
array2[3855]=30'd480046615;
array2[3856]=30'd475850257;
array2[3857]=30'd480046615;
array2[3858]=30'd475850257;
array2[3859]=30'd475850257;
array2[3860]=30'd475850257;
array2[3861]=30'd480046615;
array2[3862]=30'd480046615;
array2[3863]=30'd480046615;
array2[3864]=30'd480046615;
array2[3865]=30'd475850257;
array2[3866]=30'd480046615;
array2[3867]=30'd480046615;
array2[3868]=30'd480046615;
array2[3869]=30'd475850257;
array2[3870]=30'd475850257;
array2[3871]=30'd480046615;
array2[3872]=30'd480046615;
array2[3873]=30'd480046615;
array2[3874]=30'd480046615;
array2[3875]=30'd475850257;
array2[3876]=30'd457992679;
array2[3877]=30'd280568333;
array2[3878]=30'd631447172;
array2[3879]=30'd737318494;
array2[3880]=30'd762499681;
array2[3881]=30'd764529268;
array2[3882]=30'd737318494;
array2[3883]=30'd737318494;
array2[3884]=30'd737318494;
array2[3885]=30'd749877860;
array2[3886]=30'd762499681;
array2[3887]=30'd749877860;
array2[3888]=30'd677571193;
array2[3889]=30'd646130287;
array2[3890]=30'd631447172;
array2[3891]=30'd672348794;
array2[3892]=30'd646130287;
array2[3893]=30'd672348794;
array2[3894]=30'd606320275;
array2[3895]=30'd407216718;
array2[3896]=30'd407216718;
array2[3897]=30'd347490866;
array2[3898]=30'd260631016;
array2[3899]=30'd339244483;
array2[3900]=30'd339244483;
array2[3901]=30'd356016571;
array2[3902]=30'd364405173;
array2[3903]=30'd364405173;
array2[3904]=30'd356016571;
array2[3905]=30'd312021416;
array2[3906]=30'd339244483;
array2[3907]=30'd339244483;
array2[3908]=30'd356016571;
array2[3909]=30'd359161273;
array2[3910]=30'd339244483;
array2[3911]=30'd339244483;
array2[3912]=30'd339244483;
array2[3913]=30'd339244483;
array2[3914]=30'd260631016;
array2[3915]=30'd207191473;
array2[3916]=30'd195647926;
array2[3917]=30'd212454818;
array2[3918]=30'd212454818;
array2[3919]=30'd227159434;
array2[3920]=30'd228212100;
array2[3921]=30'd425297329;
array2[3922]=30'd338288022;
array2[3923]=30'd227165569;
array2[3924]=30'd231364996;
array2[3925]=30'd231362949;
array2[3926]=30'd301610387;
array2[3927]=30'd425297329;
array2[3928]=30'd248105365;
array2[3929]=30'd227159434;
array2[3930]=30'd234504581;
array2[3931]=30'd227165569;
array2[3932]=30'd231364996;
array2[3933]=30'd231359873;
array2[3934]=30'd230317442;
array2[3935]=30'd230317442;
array2[3936]=30'd387723742;
array2[3937]=30'd439121402;
array2[3938]=30'd439121402;
array2[3939]=30'd480046615;
array2[3940]=30'd475850257;
array2[3941]=30'd480046615;
array2[3942]=30'd475850257;
array2[3943]=30'd480046615;
array2[3944]=30'd475850257;
array2[3945]=30'd480046615;
array2[3946]=30'd480046615;
array2[3947]=30'd480046615;
array2[3948]=30'd475850257;
array2[3949]=30'd473746934;
array2[3950]=30'd439121402;
array2[3951]=30'd439121402;
array2[3952]=30'd439121402;
array2[3953]=30'd439121402;
array2[3954]=30'd439121402;
array2[3955]=30'd439121402;
array2[3956]=30'd439121402;
array2[3957]=30'd439121402;
array2[3958]=30'd439121402;
array2[3959]=30'd439121402;
array2[3960]=30'd439121402;
array2[3961]=30'd439121402;
array2[3962]=30'd475850257;
array2[3963]=30'd480046615;
array2[3964]=30'd480046615;
array2[3965]=30'd475850257;
array2[3966]=30'd475850257;
array2[3967]=30'd480046615;
array2[3968]=30'd480046615;
array2[3969]=30'd480046615;
array2[3970]=30'd480046615;
array2[3971]=30'd475850257;
array2[3972]=30'd457992679;
array2[3973]=30'd280568333;
array2[3974]=30'd646130287;
array2[3975]=30'd727851632;
array2[3976]=30'd727851632;
array2[3977]=30'd762499681;
array2[3978]=30'd749877860;
array2[3979]=30'd749877860;
array2[3980]=30'd762499681;
array2[3981]=30'd749877860;
array2[3982]=30'd762499681;
array2[3983]=30'd678602388;
array2[3984]=30'd631447172;
array2[3985]=30'd646130287;
array2[3986]=30'd565444213;
array2[3987]=30'd347490866;
array2[3988]=30'd319215128;
array2[3989]=30'd319215128;
array2[3990]=30'd319215128;
array2[3991]=30'd207191473;
array2[3992]=30'd212454818;
array2[3993]=30'd212454818;
array2[3994]=30'd254365107;
array2[3995]=30'd339244483;
array2[3996]=30'd356016571;
array2[3997]=30'd359161273;
array2[3998]=30'd356016571;
array2[3999]=30'd359161273;
array2[4000]=30'd356016571;
array2[4001]=30'd295249323;
array2[4002]=30'd339244483;
array2[4003]=30'd356016571;
array2[4004]=30'd356016571;
array2[4005]=30'd356016571;
array2[4006]=30'd339244483;
array2[4007]=30'd339244483;
array2[4008]=30'd339244483;
array2[4009]=30'd267996623;
array2[4010]=30'd228181405;
array2[4011]=30'd221916546;
array2[4012]=30'd227165569;
array2[4013]=30'd231362949;
array2[4014]=30'd256519562;
array2[4015]=30'd338288022;
array2[4016]=30'd472496545;
array2[4017]=30'd256519562;
array2[4018]=30'd228216193;
array2[4019]=30'd231359873;
array2[4020]=30'd228216193;
array2[4021]=30'd230317442;
array2[4022]=30'd230317442;
array2[4023]=30'd272255371;
array2[4024]=30'd464076202;
array2[4025]=30'd338288022;
array2[4026]=30'd228212100;
array2[4027]=30'd231362949;
array2[4028]=30'd229266819;
array2[4029]=30'd231364996;
array2[4030]=30'd229266819;
array2[4031]=30'd230317442;
array2[4032]=30'd212454818;
array2[4033]=30'd231362949;
array2[4034]=30'd307963313;
array2[4035]=30'd387723742;
array2[4036]=30'd387723742;
array2[4037]=30'd387723742;
array2[4038]=30'd387723742;
array2[4039]=30'd387723742;
array2[4040]=30'd387723742;
array2[4041]=30'd387723742;
array2[4042]=30'd387723742;
array2[4043]=30'd387723742;
array2[4044]=30'd340509129;
array2[4045]=30'd362496490;
array2[4046]=30'd232422779;
array2[4047]=30'd234504581;
array2[4048]=30'd231362949;
array2[4049]=30'd231362949;
array2[4050]=30'd229270912;
array2[4051]=30'd232417668;
array2[4052]=30'd231364996;
array2[4053]=30'd231364996;
array2[4054]=30'd234504581;
array2[4055]=30'd227165569;
array2[4056]=30'd230307208;
array2[4057]=30'd265985428;
array2[4058]=30'd387723742;
array2[4059]=30'd387723742;
array2[4060]=30'd387723742;
array2[4061]=30'd387723742;
array2[4062]=30'd387723742;
array2[4063]=30'd387723742;
array2[4064]=30'd387723742;
array2[4065]=30'd387723742;
array2[4066]=30'd387723742;
array2[4067]=30'd387723742;
array2[4068]=30'd302686639;
array2[4069]=30'd347490866;
array2[4070]=30'd646130287;
array2[4071]=30'd729975381;
array2[4072]=30'd729975381;
array2[4073]=30'd729975381;
array2[4074]=30'd737318494;
array2[4075]=30'd737318494;
array2[4076]=30'd737318494;
array2[4077]=30'd737318494;
array2[4078]=30'd677571193;
array2[4079]=30'd565444213;
array2[4080]=30'd401997362;
array2[4081]=30'd281508345;
array2[4082]=30'd281508345;
array2[4083]=30'd228181405;
array2[4084]=30'd213516691;
array2[4085]=30'd213516691;
array2[4086]=30'd213516691;
array2[4087]=30'd225072515;
array2[4088]=30'd230317442;
array2[4089]=30'd229266819;
array2[4090]=30'd234499470;
array2[4091]=30'd295249323;
array2[4092]=30'd339244483;
array2[4093]=30'd356016571;
array2[4094]=30'd356016571;
array2[4095]=30'd356016571;
array2[4096]=30'd356016571;
array2[4097]=30'd312021416;
array2[4098]=30'd295249323;
array2[4099]=30'd295249323;
array2[4100]=30'd295249323;
array2[4101]=30'd295249323;
array2[4102]=30'd248105365;
array2[4103]=30'd228181405;
array2[4104]=30'd210373000;
array2[4105]=30'd232392085;
array2[4106]=30'd232392085;
array2[4107]=30'd228216193;
array2[4108]=30'd229266819;
array2[4109]=30'd230317442;
array2[4110]=30'd256519562;
array2[4111]=30'd338288022;
array2[4112]=30'd603537847;
array2[4113]=30'd338288022;
array2[4114]=30'd221916546;
array2[4115]=30'd229270912;
array2[4116]=30'd229266819;
array2[4117]=30'd231364996;
array2[4118]=30'd229266819;
array2[4119]=30'd256519562;
array2[4120]=30'd603537847;
array2[4121]=30'd425297329;
array2[4122]=30'd227165569;
array2[4123]=30'd231362949;
array2[4124]=30'd231362949;
array2[4125]=30'd229266819;
array2[4126]=30'd231362949;
array2[4127]=30'd231362949;
array2[4128]=30'd212454818;
array2[4129]=30'd234504581;
array2[4130]=30'd227165569;
array2[4131]=30'd228216193;
array2[4132]=30'd231362949;
array2[4133]=30'd230317442;
array2[4134]=30'd231359873;
array2[4135]=30'd231362949;
array2[4136]=30'd231359873;
array2[4137]=30'd230317442;
array2[4138]=30'd231362949;
array2[4139]=30'd231362949;
array2[4140]=30'd228216193;
array2[4141]=30'd229266819;
array2[4142]=30'd231359873;
array2[4143]=30'd231364996;
array2[4144]=30'd227165569;
array2[4145]=30'd234504581;
array2[4146]=30'd231362949;
array2[4147]=30'd231362949;
array2[4148]=30'd231362949;
array2[4149]=30'd231362949;
array2[4150]=30'd231362949;
array2[4151]=30'd231362949;
array2[4152]=30'd234504581;
array2[4153]=30'd231362949;
array2[4154]=30'd231362949;
array2[4155]=30'd228212100;
array2[4156]=30'd234504581;
array2[4157]=30'd231364996;
array2[4158]=30'd227165569;
array2[4159]=30'd227165569;
array2[4160]=30'd227159434;
array2[4161]=30'd231359873;
array2[4162]=30'd213516691;
array2[4163]=30'd190356956;
array2[4164]=30'd383147560;
array2[4165]=30'd506770009;
array2[4166]=30'd631447172;
array2[4167]=30'd678604396;
array2[4168]=30'd708987491;
array2[4169]=30'd708987491;
array2[4170]=30'd729975381;
array2[4171]=30'd729975381;
array2[4172]=30'd708987491;
array2[4173]=30'd645112409;
array2[4174]=30'd506770009;
array2[4175]=30'd190356956;
array2[4176]=30'd212454818;
array2[4177]=30'd227159434;
array2[4178]=30'd231362949;
array2[4179]=30'd229266819;
array2[4180]=30'd230317442;
array2[4181]=30'd231364996;
array2[4182]=30'd231362949;
array2[4183]=30'd228216193;
array2[4184]=30'd231362949;
array2[4185]=30'd229266819;
array2[4186]=30'd228216193;
array2[4187]=30'd248105365;
array2[4188]=30'd339244483;
array2[4189]=30'd356016571;
array2[4190]=30'd359161273;
array2[4191]=30'd356016571;
array2[4192]=30'd356016571;
array2[4193]=30'd312021416;
array2[4194]=30'd295249323;
array2[4195]=30'd339244483;
array2[4196]=30'd295249323;
array2[4197]=30'd228181405;
array2[4198]=30'd228216193;
array2[4199]=30'd231359873;
array2[4200]=30'd229266819;
array2[4201]=30'd231364996;
array2[4202]=30'd231362949;
array2[4203]=30'd231362949;
array2[4204]=30'd231359873;
array2[4205]=30'd229266819;
array2[4206]=30'd230317442;
array2[4207]=30'd229266819;
array2[4208]=30'd230317442;
array2[4209]=30'd401193372;
array2[4210]=30'd338288022;
array2[4211]=30'd227165569;
array2[4212]=30'd228216193;
array2[4213]=30'd230317442;
array2[4214]=30'd272255371;
array2[4215]=30'd425297329;
array2[4216]=30'd238691720;
array2[4217]=30'd228216193;
array2[4218]=30'd231362949;
array2[4219]=30'd230317442;
array2[4220]=30'd231362949;
array2[4221]=30'd230317442;
array2[4222]=30'd231362949;
array2[4223]=30'd231362949;
array2[4224]=30'd212454818;
array2[4225]=30'd231362949;
array2[4226]=30'd231362949;
array2[4227]=30'd229266819;
array2[4228]=30'd230317442;
array2[4229]=30'd230317442;
array2[4230]=30'd231362949;
array2[4231]=30'd231364996;
array2[4232]=30'd229266819;
array2[4233]=30'd230317442;
array2[4234]=30'd231362949;
array2[4235]=30'd231364996;
array2[4236]=30'd229266819;
array2[4237]=30'd229270912;
array2[4238]=30'd227165569;
array2[4239]=30'd231362949;
array2[4240]=30'd229266819;
array2[4241]=30'd229266819;
array2[4242]=30'd229266819;
array2[4243]=30'd231364996;
array2[4244]=30'd231362949;
array2[4245]=30'd231362949;
array2[4246]=30'd231362949;
array2[4247]=30'd229266819;
array2[4248]=30'd229266819;
array2[4249]=30'd229266819;
array2[4250]=30'd231362949;
array2[4251]=30'd231359873;
array2[4252]=30'd231362949;
array2[4253]=30'd231362949;
array2[4254]=30'd231364996;
array2[4255]=30'd231362949;
array2[4256]=30'd231362949;
array2[4257]=30'd227165569;
array2[4258]=30'd207191473;
array2[4259]=30'd319215128;
array2[4260]=30'd566515308;
array2[4261]=30'd678604396;
array2[4262]=30'd538207812;
array2[4263]=30'd506770009;
array2[4264]=30'd645112409;
array2[4265]=30'd646130287;
array2[4266]=30'd678604396;
array2[4267]=30'd538207812;
array2[4268]=30'd450208341;
array2[4269]=30'd195647926;
array2[4270]=30'd207191473;
array2[4271]=30'd228212100;
array2[4272]=30'd228212100;
array2[4273]=30'd230317442;
array2[4274]=30'd231362949;
array2[4275]=30'd229266819;
array2[4276]=30'd228216193;
array2[4277]=30'd231362949;
array2[4278]=30'd231362949;
array2[4279]=30'd227165569;
array2[4280]=30'd229266819;
array2[4281]=30'd229266819;
array2[4282]=30'd231362949;
array2[4283]=30'd225072515;
array2[4284]=30'd254365107;
array2[4285]=30'd339244483;
array2[4286]=30'd356016571;
array2[4287]=30'd356016571;
array2[4288]=30'd339244483;
array2[4289]=30'd339244483;
array2[4290]=30'd254365107;
array2[4291]=30'd295249323;
array2[4292]=30'd295249323;
array2[4293]=30'd248105365;
array2[4294]=30'd232392085;
array2[4295]=30'd228216193;
array2[4296]=30'd230317442;
array2[4297]=30'd231362949;
array2[4298]=30'd231362949;
array2[4299]=30'd231362949;
array2[4300]=30'd231362949;
array2[4301]=30'd229266819;
array2[4302]=30'd229266819;
array2[4303]=30'd231362949;
array2[4304]=30'd229266819;
array2[4305]=30'd489282972;
array2[4306]=30'd464076202;
array2[4307]=30'd262793620;
array2[4308]=30'd472496545;
array2[4309]=30'd338288022;
array2[4310]=30'd338288022;
array2[4311]=30'd553231776;
array2[4312]=30'd262793620;
array2[4313]=30'd230307208;
array2[4314]=30'd234504581;
array2[4315]=30'd228216193;
array2[4316]=30'd230317442;
array2[4317]=30'd229266819;
array2[4318]=30'd231362949;
array2[4319]=30'd228212100;
array2[4320]=30'd212454818;
array2[4321]=30'd234504581;
array2[4322]=30'd231359873;
array2[4323]=30'd228216193;
array2[4324]=30'd231364996;
array2[4325]=30'd230317442;
array2[4326]=30'd229266819;
array2[4327]=30'd231362949;
array2[4328]=30'd229266819;
array2[4329]=30'd230317442;
array2[4330]=30'd231362949;
array2[4331]=30'd231362949;
array2[4332]=30'd230317442;
array2[4333]=30'd227165569;
array2[4334]=30'd234504581;
array2[4335]=30'd231362949;
array2[4336]=30'd229266819;
array2[4337]=30'd229266819;
array2[4338]=30'd230317442;
array2[4339]=30'd228216193;
array2[4340]=30'd229266819;
array2[4341]=30'd231362949;
array2[4342]=30'd230317442;
array2[4343]=30'd229266819;
array2[4344]=30'd231362949;
array2[4345]=30'd231362949;
array2[4346]=30'd231359873;
array2[4347]=30'd231362949;
array2[4348]=30'd231362949;
array2[4349]=30'd231364996;
array2[4350]=30'd231362949;
array2[4351]=30'd231362949;
array2[4352]=30'd231364996;
array2[4353]=30'd232392085;
array2[4354]=30'd190356956;
array2[4355]=30'd450208341;
array2[4356]=30'd565444213;
array2[4357]=30'd506770009;
array2[4358]=30'd260631016;
array2[4359]=30'd179916222;
array2[4360]=30'd407216718;
array2[4361]=30'd444954173;
array2[4362]=30'd444954173;
array2[4363]=30'd260631016;
array2[4364]=30'd186252693;
array2[4365]=30'd220861839;
array2[4366]=30'd229266819;
array2[4367]=30'd229266819;
array2[4368]=30'd229266819;
array2[4369]=30'd229266819;
array2[4370]=30'd231359873;
array2[4371]=30'd229266819;
array2[4372]=30'd228212100;
array2[4373]=30'd231362949;
array2[4374]=30'd229266819;
array2[4375]=30'd231362949;
array2[4376]=30'd231364996;
array2[4377]=30'd231362949;
array2[4378]=30'd234504581;
array2[4379]=30'd231362949;
array2[4380]=30'd227159434;
array2[4381]=30'd295249323;
array2[4382]=30'd356016571;
array2[4383]=30'd356016571;
array2[4384]=30'd356016571;
array2[4385]=30'd359161273;
array2[4386]=30'd295249323;
array2[4387]=30'd312021416;
array2[4388]=30'd339244483;
array2[4389]=30'd295249323;
array2[4390]=30'd228181405;
array2[4391]=30'd228216193;
array2[4392]=30'd229266819;
array2[4393]=30'd231364996;
array2[4394]=30'd231362949;
array2[4395]=30'd228216193;
array2[4396]=30'd234504581;
array2[4397]=30'd229266819;
array2[4398]=30'd229266819;
array2[4399]=30'd229266819;
array2[4400]=30'd229266819;
array2[4401]=30'd231362949;
array2[4402]=30'd227165569;
array2[4403]=30'd272255371;
array2[4404]=30'd655981997;
array2[4405]=30'd425297329;
array2[4406]=30'd228212100;
array2[4407]=30'd228212100;
array2[4408]=30'd231362949;
array2[4409]=30'd227159434;
array2[4410]=30'd228216193;
array2[4411]=30'd234504581;
array2[4412]=30'd228216193;
array2[4413]=30'd229266819;
array2[4414]=30'd229266819;
array2[4415]=30'd229266819;
array2[4416]=30'd212454818;
array2[4417]=30'd231362949;
array2[4418]=30'd231362949;
array2[4419]=30'd229266819;
array2[4420]=30'd230317442;
array2[4421]=30'd231364996;
array2[4422]=30'd228216193;
array2[4423]=30'd229266819;
array2[4424]=30'd231362949;
array2[4425]=30'd231364996;
array2[4426]=30'd231362949;
array2[4427]=30'd234504581;
array2[4428]=30'd229266819;
array2[4429]=30'd234504581;
array2[4430]=30'd231362949;
array2[4431]=30'd231362949;
array2[4432]=30'd231362949;
array2[4433]=30'd229266819;
array2[4434]=30'd231362949;
array2[4435]=30'd231364996;
array2[4436]=30'd231362949;
array2[4437]=30'd229266819;
array2[4438]=30'd231364996;
array2[4439]=30'd229266819;
array2[4440]=30'd231362949;
array2[4441]=30'd231362949;
array2[4442]=30'd229266819;
array2[4443]=30'd230317442;
array2[4444]=30'd229266819;
array2[4445]=30'd230317442;
array2[4446]=30'd231362949;
array2[4447]=30'd231362949;
array2[4448]=30'd234504581;
array2[4449]=30'd220861839;
array2[4450]=30'd281508345;
array2[4451]=30'd506770009;
array2[4452]=30'd483727963;
array2[4453]=30'd260631016;
array2[4454]=30'd228212100;
array2[4455]=30'd227165569;
array2[4456]=30'd186252693;
array2[4457]=30'd193577377;
array2[4458]=30'd212454818;
array2[4459]=30'd232392085;
array2[4460]=30'd231362949;
array2[4461]=30'd230317442;
array2[4462]=30'd231362949;
array2[4463]=30'd231362949;
array2[4464]=30'd229266819;
array2[4465]=30'd231362949;
array2[4466]=30'd230317442;
array2[4467]=30'd231362949;
array2[4468]=30'd231359873;
array2[4469]=30'd231362949;
array2[4470]=30'd231362949;
array2[4471]=30'd231364996;
array2[4472]=30'd230317442;
array2[4473]=30'd231362949;
array2[4474]=30'd231362949;
array2[4475]=30'd231362949;
array2[4476]=30'd228216193;
array2[4477]=30'd257539480;
array2[4478]=30'd312021416;
array2[4479]=30'd356016571;
array2[4480]=30'd356016571;
array2[4481]=30'd359161273;
array2[4482]=30'd312021416;
array2[4483]=30'd295249323;
array2[4484]=30'd312021416;
array2[4485]=30'd295249323;
array2[4486]=30'd228181405;
array2[4487]=30'd227159434;
array2[4488]=30'd230307208;
array2[4489]=30'd231364996;
array2[4490]=30'd230317442;
array2[4491]=30'd229266819;
array2[4492]=30'd228216193;
array2[4493]=30'd229266819;
array2[4494]=30'd229266819;
array2[4495]=30'd229266819;
array2[4496]=30'd229266819;
array2[4497]=30'd230317442;
array2[4498]=30'd231362949;
array2[4499]=30'd231359873;
array2[4500]=30'd234504581;
array2[4501]=30'd230307208;
array2[4502]=30'd228216193;
array2[4503]=30'd231362949;
array2[4504]=30'd231362949;
array2[4505]=30'd231362949;
array2[4506]=30'd231362949;
array2[4507]=30'd231364996;
array2[4508]=30'd231364996;
array2[4509]=30'd234504581;
array2[4510]=30'd231362949;
array2[4511]=30'd231362949;
array2[4512]=30'd213516691;
array2[4513]=30'd231362949;
array2[4514]=30'd231364996;
array2[4515]=30'd229266819;
array2[4516]=30'd230317442;
array2[4517]=30'd231364996;
array2[4518]=30'd229266819;
array2[4519]=30'd231362949;
array2[4520]=30'd231362949;
array2[4521]=30'd231362949;
array2[4522]=30'd231362949;
array2[4523]=30'd231362949;
array2[4524]=30'd229266819;
array2[4525]=30'd229266819;
array2[4526]=30'd230317442;
array2[4527]=30'd231364996;
array2[4528]=30'd234504581;
array2[4529]=30'd231362949;
array2[4530]=30'd234504581;
array2[4531]=30'd229266819;
array2[4532]=30'd231362949;
array2[4533]=30'd229266819;
array2[4534]=30'd231364996;
array2[4535]=30'd230317442;
array2[4536]=30'd231362949;
array2[4537]=30'd231364996;
array2[4538]=30'd229266819;
array2[4539]=30'd229266819;
array2[4540]=30'd229266819;
array2[4541]=30'd229266819;
array2[4542]=30'd229266819;
array2[4543]=30'd231359873;
array2[4544]=30'd229266819;
array2[4545]=30'd220861839;
array2[4546]=30'd281508345;
array2[4547]=30'd483727963;
array2[4548]=30'd347490866;
array2[4549]=30'd213516691;
array2[4550]=30'd230317442;
array2[4551]=30'd230317442;
array2[4552]=30'd230317442;
array2[4553]=30'd227165569;
array2[4554]=30'd230317442;
array2[4555]=30'd231359873;
array2[4556]=30'd230317442;
array2[4557]=30'd229266819;
array2[4558]=30'd231362949;
array2[4559]=30'd230317442;
array2[4560]=30'd228216193;
array2[4561]=30'd229266819;
array2[4562]=30'd231359873;
array2[4563]=30'd231364996;
array2[4564]=30'd234504581;
array2[4565]=30'd231362949;
array2[4566]=30'd231364996;
array2[4567]=30'd231362949;
array2[4568]=30'd231364996;
array2[4569]=30'd231364996;
array2[4570]=30'd230317442;
array2[4571]=30'd230317442;
array2[4572]=30'd231362949;
array2[4573]=30'd231362949;
array2[4574]=30'd248105365;
array2[4575]=30'd339244483;
array2[4576]=30'd356016571;
array2[4577]=30'd356016571;
array2[4578]=30'd295249323;
array2[4579]=30'd295249323;
array2[4580]=30'd312021416;
array2[4581]=30'd295249323;
array2[4582]=30'd254365107;
array2[4583]=30'd221916546;
array2[4584]=30'd227165569;
array2[4585]=30'd228216193;
array2[4586]=30'd230317442;
array2[4587]=30'd229266819;
array2[4588]=30'd231362949;
array2[4589]=30'd231362949;
array2[4590]=30'd230317442;
array2[4591]=30'd231362949;
array2[4592]=30'd231362949;
array2[4593]=30'd231362949;
array2[4594]=30'd229266819;
array2[4595]=30'd231362949;
array2[4596]=30'd229266819;
array2[4597]=30'd231362949;
array2[4598]=30'd231362949;
array2[4599]=30'd231362949;
array2[4600]=30'd231362949;
array2[4601]=30'd231362949;
array2[4602]=30'd231362949;
array2[4603]=30'd229266819;
array2[4604]=30'd231364996;
array2[4605]=30'd229266819;
array2[4606]=30'd230317442;
array2[4607]=30'd231364996;
array2[4608]=30'd212454818;
array2[4609]=30'd234504581;
array2[4610]=30'd231359873;
array2[4611]=30'd228216193;
array2[4612]=30'd231362949;
array2[4613]=30'd230317442;
array2[4614]=30'd231359873;
array2[4615]=30'd231362949;
array2[4616]=30'd231359873;
array2[4617]=30'd229266819;
array2[4618]=30'd231362949;
array2[4619]=30'd231362949;
array2[4620]=30'd230317442;
array2[4621]=30'd234515845;
array2[4622]=30'd227165569;
array2[4623]=30'd229266819;
array2[4624]=30'd231364996;
array2[4625]=30'd231362949;
array2[4626]=30'd231362949;
array2[4627]=30'd231362949;
array2[4628]=30'd231359873;
array2[4629]=30'd229266819;
array2[4630]=30'd229266819;
array2[4631]=30'd230317442;
array2[4632]=30'd231362949;
array2[4633]=30'd231362949;
array2[4634]=30'd229266819;
array2[4635]=30'd234504581;
array2[4636]=30'd231364996;
array2[4637]=30'd234504581;
array2[4638]=30'd229266819;
array2[4639]=30'd229266819;
array2[4640]=30'd230317442;
array2[4641]=30'd220861839;
array2[4642]=30'd190356956;
array2[4643]=30'd319215128;
array2[4644]=30'd254365107;
array2[4645]=30'd227159434;
array2[4646]=30'd231362949;
array2[4647]=30'd229266819;
array2[4648]=30'd229266819;
array2[4649]=30'd225072515;
array2[4650]=30'd228216193;
array2[4651]=30'd229266819;
array2[4652]=30'd231364996;
array2[4653]=30'd230317442;
array2[4654]=30'd228216193;
array2[4655]=30'd231362949;
array2[4656]=30'd231362949;
array2[4657]=30'd229266819;
array2[4658]=30'd229266819;
array2[4659]=30'd230317442;
array2[4660]=30'd229266819;
array2[4661]=30'd231362949;
array2[4662]=30'd231362949;
array2[4663]=30'd234504581;
array2[4664]=30'd231364996;
array2[4665]=30'd234504581;
array2[4666]=30'd231364996;
array2[4667]=30'd231364996;
array2[4668]=30'd230317442;
array2[4669]=30'd231364996;
array2[4670]=30'd238691720;
array2[4671]=30'd295249323;
array2[4672]=30'd339244483;
array2[4673]=30'd356016571;
array2[4674]=30'd339244483;
array2[4675]=30'd254365107;
array2[4676]=30'd228181405;
array2[4677]=30'd295249323;
array2[4678]=30'd267996623;
array2[4679]=30'd228181405;
array2[4680]=30'd221916546;
array2[4681]=30'd228212100;
array2[4682]=30'd231364996;
array2[4683]=30'd228216193;
array2[4684]=30'd230317442;
array2[4685]=30'd231362949;
array2[4686]=30'd231362949;
array2[4687]=30'd225072515;
array2[4688]=30'd231362949;
array2[4689]=30'd231362949;
array2[4690]=30'd234504581;
array2[4691]=30'd229266819;
array2[4692]=30'd230317442;
array2[4693]=30'd229266819;
array2[4694]=30'd231362949;
array2[4695]=30'd231362949;
array2[4696]=30'd231362949;
array2[4697]=30'd234504581;
array2[4698]=30'd231362949;
array2[4699]=30'd231364996;
array2[4700]=30'd231362949;
array2[4701]=30'd231364996;
array2[4702]=30'd231362949;
array2[4703]=30'd231364996;
array2[4704]=30'd212454818;
array2[4705]=30'd234504581;
array2[4706]=30'd227165569;
array2[4707]=30'd228216193;
array2[4708]=30'd231362949;
array2[4709]=30'd230317442;
array2[4710]=30'd231359873;
array2[4711]=30'd231362949;
array2[4712]=30'd231359873;
array2[4713]=30'd230317442;
array2[4714]=30'd231362949;
array2[4715]=30'd231362949;
array2[4716]=30'd230317442;
array2[4717]=30'd234515845;
array2[4718]=30'd228212100;
array2[4719]=30'd231359873;
array2[4720]=30'd231364996;
array2[4721]=30'd231362949;
array2[4722]=30'd231362949;
array2[4723]=30'd231362949;
array2[4724]=30'd231359873;
array2[4725]=30'd231362949;
array2[4726]=30'd231362949;
array2[4727]=30'd230317442;
array2[4728]=30'd231364996;
array2[4729]=30'd231362949;
array2[4730]=30'd234504581;
array2[4731]=30'd231362949;
array2[4732]=30'd229266819;
array2[4733]=30'd234504581;
array2[4734]=30'd229266819;
array2[4735]=30'd231362949;
array2[4736]=30'd231364996;
array2[4737]=30'd221916546;
array2[4738]=30'd179916222;
array2[4739]=30'd249001484;
array2[4740]=30'd193577377;
array2[4741]=30'd228212100;
array2[4742]=30'd231362949;
array2[4743]=30'd234504581;
array2[4744]=30'd229266819;
array2[4745]=30'd229266819;
array2[4746]=30'd231362949;
array2[4747]=30'd231362949;
array2[4748]=30'd231362949;
array2[4749]=30'd231364996;
array2[4750]=30'd230317442;
array2[4751]=30'd234504581;
array2[4752]=30'd231359873;
array2[4753]=30'd231362949;
array2[4754]=30'd231362949;
array2[4755]=30'd231362949;
array2[4756]=30'd231362949;
array2[4757]=30'd231362949;
array2[4758]=30'd231362949;
array2[4759]=30'd231362949;
array2[4760]=30'd231362949;
array2[4761]=30'd229266819;
array2[4762]=30'd229266819;
array2[4763]=30'd231364996;
array2[4764]=30'd231362949;
array2[4765]=30'd231364996;
array2[4766]=30'd231362949;
array2[4767]=30'd240774546;
array2[4768]=30'd295249323;
array2[4769]=30'd339244483;
array2[4770]=30'd295249323;
array2[4771]=30'd228181405;
array2[4772]=30'd230307208;
array2[4773]=30'd248105365;
array2[4774]=30'd248105365;
array2[4775]=30'd240774546;
array2[4776]=30'd221916546;
array2[4777]=30'd231362949;
array2[4778]=30'd229266819;
array2[4779]=30'd230317442;
array2[4780]=30'd231362949;
array2[4781]=30'd228212100;
array2[4782]=30'd231362949;
array2[4783]=30'd228216193;
array2[4784]=30'd231362949;
array2[4785]=30'd231362949;
array2[4786]=30'd231364996;
array2[4787]=30'd230317442;
array2[4788]=30'd234504581;
array2[4789]=30'd234504581;
array2[4790]=30'd231362949;
array2[4791]=30'd231362949;
array2[4792]=30'd234504581;
array2[4793]=30'd231362949;
array2[4794]=30'd231362949;
array2[4795]=30'd229266819;
array2[4796]=30'd231362949;
array2[4797]=30'd234504581;
array2[4798]=30'd231362949;
array2[4799]=30'd234504581;
array2[4800]=30'd212454818;
array2[4801]=30'd234504581;
array2[4802]=30'd231359873;
array2[4803]=30'd228216193;
array2[4804]=30'd231362949;
array2[4805]=30'd230317442;
array2[4806]=30'd229266819;
array2[4807]=30'd231362949;
array2[4808]=30'd231362949;
array2[4809]=30'd231364996;
array2[4810]=30'd231362949;
array2[4811]=30'd231362949;
array2[4812]=30'd230317442;
array2[4813]=30'd229270912;
array2[4814]=30'd228216193;
array2[4815]=30'd229266819;
array2[4816]=30'd231364996;
array2[4817]=30'd231362949;
array2[4818]=30'd228216193;
array2[4819]=30'd229266819;
array2[4820]=30'd231362949;
array2[4821]=30'd229266819;
array2[4822]=30'd229266819;
array2[4823]=30'd230317442;
array2[4824]=30'd231362949;
array2[4825]=30'd231362949;
array2[4826]=30'd234504581;
array2[4827]=30'd231362949;
array2[4828]=30'd231362949;
array2[4829]=30'd231362949;
array2[4830]=30'd231362949;
array2[4831]=30'd231364996;
array2[4832]=30'd231362949;
array2[4833]=30'd231362949;
array2[4834]=30'd220861839;
array2[4835]=30'd195647926;
array2[4836]=30'd213516691;
array2[4837]=30'd228216193;
array2[4838]=30'd231362949;
array2[4839]=30'd231364996;
array2[4840]=30'd228216193;
array2[4841]=30'd231362949;
array2[4842]=30'd230307208;
array2[4843]=30'd229266819;
array2[4844]=30'd229266819;
array2[4845]=30'd229266819;
array2[4846]=30'd229266819;
array2[4847]=30'd231364996;
array2[4848]=30'd231362949;
array2[4849]=30'd234504581;
array2[4850]=30'd231362949;
array2[4851]=30'd234504581;
array2[4852]=30'd231362949;
array2[4853]=30'd230317442;
array2[4854]=30'd231362949;
array2[4855]=30'd229266819;
array2[4856]=30'd231364996;
array2[4857]=30'd231362949;
array2[4858]=30'd231364996;
array2[4859]=30'd231364996;
array2[4860]=30'd231362949;
array2[4861]=30'd231364996;
array2[4862]=30'd231364996;
array2[4863]=30'd229266819;
array2[4864]=30'd227159434;
array2[4865]=30'd227159434;
array2[4866]=30'd257539480;
array2[4867]=30'd232392085;
array2[4868]=30'd228216193;
array2[4869]=30'd230307208;
array2[4870]=30'd228216193;
array2[4871]=30'd231362949;
array2[4872]=30'd229266819;
array2[4873]=30'd231364996;
array2[4874]=30'd230317442;
array2[4875]=30'd231362949;
array2[4876]=30'd231362949;
array2[4877]=30'd228216193;
array2[4878]=30'd229266819;
array2[4879]=30'd229266819;
array2[4880]=30'd229266819;
array2[4881]=30'd231362949;
array2[4882]=30'd231362949;
array2[4883]=30'd231362949;
array2[4884]=30'd234504581;
array2[4885]=30'd231362949;
array2[4886]=30'd234504581;
array2[4887]=30'd231364996;
array2[4888]=30'd231364996;
array2[4889]=30'd229266819;
array2[4890]=30'd230317442;
array2[4891]=30'd231364996;
array2[4892]=30'd229266819;
array2[4893]=30'd231364996;
array2[4894]=30'd231362949;
array2[4895]=30'd231362949;
array2[4896]=30'd212454818;
array2[4897]=30'd234504581;
array2[4898]=30'd231362949;
array2[4899]=30'd228216193;
array2[4900]=30'd229266819;
array2[4901]=30'd230317442;
array2[4902]=30'd228216193;
array2[4903]=30'd229266819;
array2[4904]=30'd229266819;
array2[4905]=30'd230317442;
array2[4906]=30'd231362949;
array2[4907]=30'd231362949;
array2[4908]=30'd230317442;
array2[4909]=30'd229270912;
array2[4910]=30'd228216193;
array2[4911]=30'd230317442;
array2[4912]=30'd229266819;
array2[4913]=30'd229266819;
array2[4914]=30'd229266819;
array2[4915]=30'd231364996;
array2[4916]=30'd231362949;
array2[4917]=30'd231362949;
array2[4918]=30'd231362949;
array2[4919]=30'd230317442;
array2[4920]=30'd229266819;
array2[4921]=30'd231362949;
array2[4922]=30'd231364996;
array2[4923]=30'd231362949;
array2[4924]=30'd229266819;
array2[4925]=30'd231359873;
array2[4926]=30'd231364996;
array2[4927]=30'd231362949;
array2[4928]=30'd231362949;
array2[4929]=30'd231364996;
array2[4930]=30'd231362949;
array2[4931]=30'd228216193;
array2[4932]=30'd231364996;
array2[4933]=30'd229266819;
array2[4934]=30'd230317442;
array2[4935]=30'd229266819;
array2[4936]=30'd231362949;
array2[4937]=30'd231362949;
array2[4938]=30'd228216193;
array2[4939]=30'd231362949;
array2[4940]=30'd231362949;
array2[4941]=30'd231364996;
array2[4942]=30'd231362949;
array2[4943]=30'd231364996;
array2[4944]=30'd231362949;
array2[4945]=30'd229266819;
array2[4946]=30'd231364996;
array2[4947]=30'd229266819;
array2[4948]=30'd230317442;
array2[4949]=30'd231362949;
array2[4950]=30'd231362949;
array2[4951]=30'd231362949;
array2[4952]=30'd231362949;
array2[4953]=30'd231362949;
array2[4954]=30'd231362949;
array2[4955]=30'd229270912;
array2[4956]=30'd231362949;
array2[4957]=30'd231362949;
array2[4958]=30'd231364996;
array2[4959]=30'd229266819;
array2[4960]=30'd230317442;
array2[4961]=30'd229266819;
array2[4962]=30'd229266819;
array2[4963]=30'd231362949;
array2[4964]=30'd231362949;
array2[4965]=30'd231362949;
array2[4966]=30'd231364996;
array2[4967]=30'd231364996;
array2[4968]=30'd231364996;
array2[4969]=30'd229270912;
array2[4970]=30'd230317442;
array2[4971]=30'd229266819;
array2[4972]=30'd231364996;
array2[4973]=30'd229266819;
array2[4974]=30'd229270912;
array2[4975]=30'd229266819;
array2[4976]=30'd229266819;
array2[4977]=30'd229266819;
array2[4978]=30'd231362949;
array2[4979]=30'd229266819;
array2[4980]=30'd231362949;
array2[4981]=30'd229266819;
array2[4982]=30'd230317442;
array2[4983]=30'd229266819;
array2[4984]=30'd231362949;
array2[4985]=30'd231364996;
array2[4986]=30'd229266819;
array2[4987]=30'd231362949;
array2[4988]=30'd229266819;
array2[4989]=30'd230317442;
array2[4990]=30'd229266819;
array2[4991]=30'd229270912;
array2[4992]=30'd212454818;
array2[4993]=30'd231362949;
array2[4994]=30'd231362949;
array2[4995]=30'd229266819;
array2[4996]=30'd230317442;
array2[4997]=30'd231364996;
array2[4998]=30'd231359873;
array2[4999]=30'd230317442;
array2[5000]=30'd231362949;
array2[5001]=30'd229266819;
array2[5002]=30'd231362949;
array2[5003]=30'd231362949;
array2[5004]=30'd231362949;
array2[5005]=30'd229270912;
array2[5006]=30'd228216193;
array2[5007]=30'd230317442;
array2[5008]=30'd231359873;
array2[5009]=30'd231362949;
array2[5010]=30'd231359873;
array2[5011]=30'd231362949;
array2[5012]=30'd231359873;
array2[5013]=30'd229266819;
array2[5014]=30'd229266819;
array2[5015]=30'd231362949;
array2[5016]=30'd231362949;
array2[5017]=30'd231362949;
array2[5018]=30'd231362949;
array2[5019]=30'd231362949;
array2[5020]=30'd231359873;
array2[5021]=30'd229266819;
array2[5022]=30'd231362949;
array2[5023]=30'd228216193;
array2[5024]=30'd229266819;
array2[5025]=30'd231362949;
array2[5026]=30'd234504581;
array2[5027]=30'd231362949;
array2[5028]=30'd231364996;
array2[5029]=30'd231364996;
array2[5030]=30'd231362949;
array2[5031]=30'd234504581;
array2[5032]=30'd231362949;
array2[5033]=30'd231362949;
array2[5034]=30'd234504581;
array2[5035]=30'd231362949;
array2[5036]=30'd231362949;
array2[5037]=30'd231362949;
array2[5038]=30'd231362949;
array2[5039]=30'd234504581;
array2[5040]=30'd231362949;
array2[5041]=30'd231362949;
array2[5042]=30'd231362949;
array2[5043]=30'd231362949;
array2[5044]=30'd231362949;
array2[5045]=30'd228216193;
array2[5046]=30'd231362949;
array2[5047]=30'd231362949;
array2[5048]=30'd231359873;
array2[5049]=30'd231362949;
array2[5050]=30'd231364996;
array2[5051]=30'd231364996;
array2[5052]=30'd231362949;
array2[5053]=30'd256519562;
array2[5054]=30'd256519562;
array2[5055]=30'd238691720;
array2[5056]=30'd231362949;
array2[5057]=30'd228216193;
array2[5058]=30'd231364996;
array2[5059]=30'd230317442;
array2[5060]=30'd231362949;
array2[5061]=30'd231362949;
array2[5062]=30'd227165569;
array2[5063]=30'd231362949;
array2[5064]=30'd231362949;
array2[5065]=30'd231362949;
array2[5066]=30'd229266819;
array2[5067]=30'd231362949;
array2[5068]=30'd229266819;
array2[5069]=30'd231362949;
array2[5070]=30'd231362949;
array2[5071]=30'd228216193;
array2[5072]=30'd231362949;
array2[5073]=30'd229266819;
array2[5074]=30'd230317442;
array2[5075]=30'd234504581;
array2[5076]=30'd231359873;
array2[5077]=30'd231362949;
array2[5078]=30'd231364996;
array2[5079]=30'd231362949;
array2[5080]=30'd234504581;
array2[5081]=30'd231362949;
array2[5082]=30'd231362949;
array2[5083]=30'd231362949;
array2[5084]=30'd231362949;
array2[5085]=30'd230317442;
array2[5086]=30'd229270912;
array2[5087]=30'd231364996;
array2[5088]=30'd213516691;
array2[5089]=30'd234504581;
array2[5090]=30'd231362949;
array2[5091]=30'd229266819;
array2[5092]=30'd231364996;
array2[5093]=30'd230317442;
array2[5094]=30'd229266819;
array2[5095]=30'd229266819;
array2[5096]=30'd229266819;
array2[5097]=30'd228212100;
array2[5098]=30'd230317442;
array2[5099]=30'd231362949;
array2[5100]=30'd230317442;
array2[5101]=30'd229270912;
array2[5102]=30'd228212100;
array2[5103]=30'd230317442;
array2[5104]=30'd230317442;
array2[5105]=30'd230317442;
array2[5106]=30'd227159434;
array2[5107]=30'd225072515;
array2[5108]=30'd229266819;
array2[5109]=30'd231364996;
array2[5110]=30'd230317442;
array2[5111]=30'd228216193;
array2[5112]=30'd231362949;
array2[5113]=30'd231359873;
array2[5114]=30'd229266819;
array2[5115]=30'd229266819;
array2[5116]=30'd229266819;
array2[5117]=30'd231362949;
array2[5118]=30'd231362949;
array2[5119]=30'd234504581;
array2[5120]=30'd234504581;
array2[5121]=30'd231364996;
array2[5122]=30'd234504581;
array2[5123]=30'd231364996;
array2[5124]=30'd231364996;
array2[5125]=30'd230317442;
array2[5126]=30'd229270912;
array2[5127]=30'd231364996;
array2[5128]=30'd229266819;
array2[5129]=30'd229270912;
array2[5130]=30'd231362949;
array2[5131]=30'd231362949;
array2[5132]=30'd231362949;
array2[5133]=30'd230317442;
array2[5134]=30'd229266819;
array2[5135]=30'd231364996;
array2[5136]=30'd230317442;
array2[5137]=30'd230307208;
array2[5138]=30'd228216193;
array2[5139]=30'd229266819;
array2[5140]=30'd230317442;
array2[5141]=30'd229266819;
array2[5142]=30'd231362949;
array2[5143]=30'd229266819;
array2[5144]=30'd231362949;
array2[5145]=30'd256519562;
array2[5146]=30'd227165569;
array2[5147]=30'd231362949;
array2[5148]=30'd229270912;
array2[5149]=30'd338288022;
array2[5150]=30'd664345022;
array2[5151]=30'd281654691;
array2[5152]=30'd234504581;
array2[5153]=30'd231359873;
array2[5154]=30'd229270912;
array2[5155]=30'd230317442;
array2[5156]=30'd229266819;
array2[5157]=30'd229270912;
array2[5158]=30'd231362949;
array2[5159]=30'd228216193;
array2[5160]=30'd234504581;
array2[5161]=30'd229266819;
array2[5162]=30'd230317442;
array2[5163]=30'd229266819;
array2[5164]=30'd229266819;
array2[5165]=30'd231362949;
array2[5166]=30'd231362949;
array2[5167]=30'd234504581;
array2[5168]=30'd231362949;
array2[5169]=30'd231362949;
array2[5170]=30'd231362949;
array2[5171]=30'd231364996;
array2[5172]=30'd229266819;
array2[5173]=30'd230317442;
array2[5174]=30'd232417668;
array2[5175]=30'd231359873;
array2[5176]=30'd230317442;
array2[5177]=30'd231364996;
array2[5178]=30'd231362949;
array2[5179]=30'd229266819;
array2[5180]=30'd231362949;
array2[5181]=30'd229266819;
array2[5182]=30'd230317442;
array2[5183]=30'd231362949;
array2[5184]=30'd193577377;
array2[5185]=30'd234504581;
array2[5186]=30'd227165569;
array2[5187]=30'd228216193;
array2[5188]=30'd228216193;
array2[5189]=30'd228216193;
array2[5190]=30'd229266819;
array2[5191]=30'd231362949;
array2[5192]=30'd234504581;
array2[5193]=30'd229266819;
array2[5194]=30'd231364996;
array2[5195]=30'd230317442;
array2[5196]=30'd231362949;
array2[5197]=30'd231362949;
array2[5198]=30'd231362949;
array2[5199]=30'd231362949;
array2[5200]=30'd231362949;
array2[5201]=30'd229266819;
array2[5202]=30'd228216193;
array2[5203]=30'd229266819;
array2[5204]=30'd229266819;
array2[5205]=30'd231359873;
array2[5206]=30'd231362949;
array2[5207]=30'd231364996;
array2[5208]=30'd230317442;
array2[5209]=30'd229266819;
array2[5210]=30'd231362949;
array2[5211]=30'd231362949;
array2[5212]=30'd231364996;
array2[5213]=30'd231362949;
array2[5214]=30'd231362949;
array2[5215]=30'd228216193;
array2[5216]=30'd231359873;
array2[5217]=30'd231362949;
array2[5218]=30'd231362949;
array2[5219]=30'd231359873;
array2[5220]=30'd231362949;
array2[5221]=30'd231364996;
array2[5222]=30'd231362949;
array2[5223]=30'd229266819;
array2[5224]=30'd234504581;
array2[5225]=30'd230317442;
array2[5226]=30'd229266819;
array2[5227]=30'd229266819;
array2[5228]=30'd231362949;
array2[5229]=30'd228216193;
array2[5230]=30'd231359873;
array2[5231]=30'd229266819;
array2[5232]=30'd231362949;
array2[5233]=30'd231362949;
array2[5234]=30'd234504581;
array2[5235]=30'd229266819;
array2[5236]=30'd229270912;
array2[5237]=30'd231364996;
array2[5238]=30'd231362949;
array2[5239]=30'd231362949;
array2[5240]=30'd230317442;
array2[5241]=30'd231362949;
array2[5242]=30'd231362949;
array2[5243]=30'd229266819;
array2[5244]=30'd227165569;
array2[5245]=30'd229266819;
array2[5246]=30'd229266819;
array2[5247]=30'd231362949;
array2[5248]=30'd231362949;
array2[5249]=30'd231362949;
array2[5250]=30'd229266819;
array2[5251]=30'd230317442;
array2[5252]=30'd231362949;
array2[5253]=30'd231362949;
array2[5254]=30'd229266819;
array2[5255]=30'd230317442;
array2[5256]=30'd231362949;
array2[5257]=30'd229266819;
array2[5258]=30'd231362949;
array2[5259]=30'd228216193;
array2[5260]=30'd229266819;
array2[5261]=30'd231362949;
array2[5262]=30'd231362949;
array2[5263]=30'd231362949;
array2[5264]=30'd272255371;
array2[5265]=30'd231362949;
array2[5266]=30'd256519562;
array2[5267]=30'd405404052;
array2[5268]=30'd272255371;
array2[5269]=30'd234504581;
array2[5270]=30'd272255371;
array2[5271]=30'd227165569;
array2[5272]=30'd229266819;
array2[5273]=30'd230317442;
array2[5274]=30'd231364996;
array2[5275]=30'd230317442;
array2[5276]=30'd231364996;
array2[5277]=30'd472496545;
array2[5278]=30'd747191732;
array2[5279]=30'd256519562;
array2[5280]=30'd193577377;
array2[5281]=30'd227165569;
array2[5282]=30'd230307208;
array2[5283]=30'd231362949;
array2[5284]=30'd229266819;
array2[5285]=30'd229266819;
array2[5286]=30'd229266819;
array2[5287]=30'd231359873;
array2[5288]=30'd229266819;
array2[5289]=30'd231362949;
array2[5290]=30'd231362949;
array2[5291]=30'd231362949;
array2[5292]=30'd228216193;
array2[5293]=30'd234504581;
array2[5294]=30'd231359873;
array2[5295]=30'd231362949;
array2[5296]=30'd231362949;
array2[5297]=30'd230317442;
array2[5298]=30'd231364996;
array2[5299]=30'd229266819;
array2[5300]=30'd227159434;
array2[5301]=30'd220861839;
array2[5302]=30'd221916546;
array2[5303]=30'd227159434;
array2[5304]=30'd227165569;
array2[5305]=30'd228216193;
array2[5306]=30'd228216193;
array2[5307]=30'd231364996;
array2[5308]=30'd231362949;
array2[5309]=30'd231362949;
array2[5310]=30'd231362949;
array2[5311]=30'd228216193;
array2[5312]=30'd231362949;
array2[5313]=30'd230317442;
array2[5314]=30'd230317442;
array2[5315]=30'd230317442;
array2[5316]=30'd229266819;
array2[5317]=30'd230317442;
array2[5318]=30'd231362949;
array2[5319]=30'd231362949;
array2[5320]=30'd231362949;
array2[5321]=30'd229266819;
array2[5322]=30'd228216193;
array2[5323]=30'd230317442;
array2[5324]=30'd229266819;
array2[5325]=30'd231362949;
array2[5326]=30'd228216193;
array2[5327]=30'd228216193;
array2[5328]=30'd229266819;
array2[5329]=30'd231362949;
array2[5330]=30'd231362949;
array2[5331]=30'd231362949;
array2[5332]=30'd230317442;
array2[5333]=30'd231362949;
array2[5334]=30'd231362949;
array2[5335]=30'd229266819;
array2[5336]=30'd229266819;
array2[5337]=30'd231362949;
array2[5338]=30'd229266819;
array2[5339]=30'd231362949;
array2[5340]=30'd229266819;
array2[5341]=30'd231362949;
array2[5342]=30'd229266819;
array2[5343]=30'd231359873;
array2[5344]=30'd231364996;
array2[5345]=30'd231362949;
array2[5346]=30'd229266819;
array2[5347]=30'd231362949;
array2[5348]=30'd231359873;
array2[5349]=30'd231362949;
array2[5350]=30'd231362949;
array2[5351]=30'd231362949;
array2[5352]=30'd231362949;
array2[5353]=30'd231362949;
array2[5354]=30'd231359873;
array2[5355]=30'd231362949;
array2[5356]=30'd231364996;
array2[5357]=30'd231362949;
array2[5358]=30'd229266819;
array2[5359]=30'd229266819;
array2[5360]=30'd229266819;
array2[5361]=30'd231359873;
array2[5362]=30'd256519562;
array2[5363]=30'd377085336;
array2[5364]=30'd256519562;
array2[5365]=30'd228216193;
array2[5366]=30'd231362949;
array2[5367]=30'd231362949;
array2[5368]=30'd231362949;
array2[5369]=30'd230317442;
array2[5370]=30'd231362949;
array2[5371]=30'd231362949;
array2[5372]=30'd229266819;
array2[5373]=30'd338288022;
array2[5374]=30'd472496545;
array2[5375]=30'd256519562;
array2[5376]=30'd193577377;
array2[5377]=30'd234504581;
array2[5378]=30'd227165569;
array2[5379]=30'd228216193;
array2[5380]=30'd229266819;
array2[5381]=30'd231362949;
array2[5382]=30'd231362949;
array2[5383]=30'd231362949;
array2[5384]=30'd229266819;
array2[5385]=30'd231362949;
array2[5386]=30'd230317442;
array2[5387]=30'd231362949;
array2[5388]=30'd229266819;
array2[5389]=30'd229266819;
array2[5390]=30'd229270912;
array2[5391]=30'd231364996;
array2[5392]=30'd229266819;
array2[5393]=30'd230317442;
array2[5394]=30'd231364996;
array2[5395]=30'd234504581;
array2[5396]=30'd179916222;
array2[5397]=30'd383147560;
array2[5398]=30'd407216718;
array2[5399]=30'd347490866;
array2[5400]=30'd193577377;
array2[5401]=30'd186252693;
array2[5402]=30'd220861839;
array2[5403]=30'd232417668;
array2[5404]=30'd228216193;
array2[5405]=30'd230317442;
array2[5406]=30'd231362949;
array2[5407]=30'd230317442;
array2[5408]=30'd231362949;
array2[5409]=30'd230317442;
array2[5410]=30'd231362949;
array2[5411]=30'd230317442;
array2[5412]=30'd229266819;
array2[5413]=30'd229270912;
array2[5414]=30'd231364996;
array2[5415]=30'd229266819;
array2[5416]=30'd231362949;
array2[5417]=30'd231362949;
array2[5418]=30'd231362949;
array2[5419]=30'd231364996;
array2[5420]=30'd231362949;
array2[5421]=30'd230317442;
array2[5422]=30'd231362949;
array2[5423]=30'd231362949;
array2[5424]=30'd231359873;
array2[5425]=30'd230317442;
array2[5426]=30'd231362949;
array2[5427]=30'd229266819;
array2[5428]=30'd231362949;
array2[5429]=30'd230317442;
array2[5430]=30'd231362949;
array2[5431]=30'd231362949;
array2[5432]=30'd231362949;
array2[5433]=30'd228216193;
array2[5434]=30'd229266819;
array2[5435]=30'd229266819;
array2[5436]=30'd229266819;
array2[5437]=30'd231362949;
array2[5438]=30'd231359873;
array2[5439]=30'd231359873;
array2[5440]=30'd229266819;
array2[5441]=30'd231362949;
array2[5442]=30'd230317442;
array2[5443]=30'd231362949;
array2[5444]=30'd231362949;
array2[5445]=30'd231362949;
array2[5446]=30'd230317442;
array2[5447]=30'd230317442;
array2[5448]=30'd231362949;
array2[5449]=30'd229266819;
array2[5450]=30'd229266819;
array2[5451]=30'd230317442;
array2[5452]=30'd229266819;
array2[5453]=30'd231364996;
array2[5454]=30'd229266819;
array2[5455]=30'd229266819;
array2[5456]=30'd231362949;
array2[5457]=30'd229266819;
array2[5458]=30'd231362949;
array2[5459]=30'd230317442;
array2[5460]=30'd231362949;
array2[5461]=30'd229266819;
array2[5462]=30'd231362949;
array2[5463]=30'd230317442;
array2[5464]=30'd231364996;
array2[5465]=30'd229266819;
array2[5466]=30'd229266819;
array2[5467]=30'd231362949;
array2[5468]=30'd228216193;
array2[5469]=30'd228216193;
array2[5470]=30'd229266819;
array2[5471]=30'd229266819;
array2[5472]=30'd193577377;
array2[5473]=30'd234504581;
array2[5474]=30'd227165569;
array2[5475]=30'd228216193;
array2[5476]=30'd230317442;
array2[5477]=30'd231364996;
array2[5478]=30'd231364996;
array2[5479]=30'd231362949;
array2[5480]=30'd229266819;
array2[5481]=30'd231362949;
array2[5482]=30'd231362949;
array2[5483]=30'd231362949;
array2[5484]=30'd230317442;
array2[5485]=30'd301610387;
array2[5486]=30'd664345022;
array2[5487]=30'd377085336;
array2[5488]=30'd227165569;
array2[5489]=30'd228216193;
array2[5490]=30'd229266819;
array2[5491]=30'd231362949;
array2[5492]=30'd179916222;
array2[5493]=30'd646130287;
array2[5494]=30'd764529268;
array2[5495]=30'd677571193;
array2[5496]=30'd483727963;
array2[5497]=30'd483727963;
array2[5498]=30'd260631016;
array2[5499]=30'd193577377;
array2[5500]=30'd193577377;
array2[5501]=30'd225072515;
array2[5502]=30'd228216193;
array2[5503]=30'd231362949;
array2[5504]=30'd231362949;
array2[5505]=30'd229266819;
array2[5506]=30'd231364996;
array2[5507]=30'd231364996;
array2[5508]=30'd256519562;
array2[5509]=30'd603537847;
array2[5510]=30'd472496545;
array2[5511]=30'd229270912;
array2[5512]=30'd231362949;
array2[5513]=30'd231362949;
array2[5514]=30'd231364996;
array2[5515]=30'd231364996;
array2[5516]=30'd231364996;
array2[5517]=30'd229266819;
array2[5518]=30'd229266819;
array2[5519]=30'd231362949;
array2[5520]=30'd229266819;
array2[5521]=30'd231362949;
array2[5522]=30'd231364996;
array2[5523]=30'd231362949;
array2[5524]=30'd230317442;
array2[5525]=30'd231362949;
array2[5526]=30'd231362949;
array2[5527]=30'd231362949;
array2[5528]=30'd229266819;
array2[5529]=30'd230317442;
array2[5530]=30'd231362949;
array2[5531]=30'd231362949;
array2[5532]=30'd231364996;
array2[5533]=30'd229266819;
array2[5534]=30'd229266819;
array2[5535]=30'd231362949;
array2[5536]=30'd231362949;
array2[5537]=30'd230317442;
array2[5538]=30'd229266819;
array2[5539]=30'd229266819;
array2[5540]=30'd231364996;
array2[5541]=30'd229266819;
array2[5542]=30'd229266819;
array2[5543]=30'd231362949;
array2[5544]=30'd229266819;
array2[5545]=30'd231362949;
array2[5546]=30'd230317442;
array2[5547]=30'd231362949;
array2[5548]=30'd228216193;
array2[5549]=30'd231362949;
array2[5550]=30'd229266819;
array2[5551]=30'd230317442;
array2[5552]=30'd231362949;
array2[5553]=30'd231364996;
array2[5554]=30'd231362949;
array2[5555]=30'd229266819;
array2[5556]=30'd231362949;
array2[5557]=30'd230317442;
array2[5558]=30'd229266819;
array2[5559]=30'd229266819;
array2[5560]=30'd230317442;
array2[5561]=30'd229266819;
array2[5562]=30'd231362949;
array2[5563]=30'd231362949;
array2[5564]=30'd230317442;
array2[5565]=30'd231362949;
array2[5566]=30'd231362949;
array2[5567]=30'd230317442;
array2[5568]=30'd193577377;
array2[5569]=30'd234504581;
array2[5570]=30'd227165569;
array2[5571]=30'd228216193;
array2[5572]=30'd230317442;
array2[5573]=30'd231362949;
array2[5574]=30'd230317442;
array2[5575]=30'd231362949;
array2[5576]=30'd228216193;
array2[5577]=30'd231362949;
array2[5578]=30'd231362949;
array2[5579]=30'd231362949;
array2[5580]=30'd229266819;
array2[5581]=30'd272255371;
array2[5582]=30'd532258209;
array2[5583]=30'd338288022;
array2[5584]=30'd227159434;
array2[5585]=30'd231364996;
array2[5586]=30'd231362949;
array2[5587]=30'd231364996;
array2[5588]=30'd179916222;
array2[5589]=30'd708987491;
array2[5590]=30'd790726247;
array2[5591]=30'd790726247;
array2[5592]=30'd790726247;
array2[5593]=30'd790726247;
array2[5594]=30'd566515308;
array2[5595]=30'd538207812;
array2[5596]=30'd483727963;
array2[5597]=30'd195647926;
array2[5598]=30'd207191473;
array2[5599]=30'd228181405;
array2[5600]=30'd230307208;
array2[5601]=30'd228216193;
array2[5602]=30'd229266819;
array2[5603]=30'd229266819;
array2[5604]=30'd256519562;
array2[5605]=30'd489282972;
array2[5606]=30'd401193372;
array2[5607]=30'd227159434;
array2[5608]=30'd228216193;
array2[5609]=30'd228216193;
array2[5610]=30'd229266819;
array2[5611]=30'd230317442;
array2[5612]=30'd231364996;
array2[5613]=30'd231362949;
array2[5614]=30'd229266819;
array2[5615]=30'd229266819;
array2[5616]=30'd229266819;
array2[5617]=30'd229266819;
array2[5618]=30'd231362949;
array2[5619]=30'd231362949;
array2[5620]=30'd229266819;
array2[5621]=30'd231364996;
array2[5622]=30'd231362949;
array2[5623]=30'd229266819;
array2[5624]=30'd231362949;
array2[5625]=30'd231364996;
array2[5626]=30'd231362949;
array2[5627]=30'd231364996;
array2[5628]=30'd231362949;
array2[5629]=30'd228216193;
array2[5630]=30'd231362949;
array2[5631]=30'd229266819;
array2[5632]=30'd231362949;
array2[5633]=30'd231362949;
array2[5634]=30'd228216193;
array2[5635]=30'd229266819;
array2[5636]=30'd234504581;
array2[5637]=30'd231362949;
array2[5638]=30'd231364996;
array2[5639]=30'd229266819;
array2[5640]=30'd228216193;
array2[5641]=30'd229266819;
array2[5642]=30'd231362949;
array2[5643]=30'd231362949;
array2[5644]=30'd231362949;
array2[5645]=30'd229266819;
array2[5646]=30'd228216193;
array2[5647]=30'd229266819;
array2[5648]=30'd229266819;
array2[5649]=30'd229266819;
array2[5650]=30'd231362949;
array2[5651]=30'd228216193;
array2[5652]=30'd231362949;
array2[5653]=30'd231362949;
array2[5654]=30'd231362949;
array2[5655]=30'd231362949;
array2[5656]=30'd231364996;
array2[5657]=30'd229270912;
array2[5658]=30'd231362949;
array2[5659]=30'd229266819;
array2[5660]=30'd231362949;
array2[5661]=30'd231362949;
array2[5662]=30'd230317442;
array2[5663]=30'd231362949;
array2[5664]=30'd193577377;
array2[5665]=30'd234504581;
array2[5666]=30'd227165569;
array2[5667]=30'd228216193;
array2[5668]=30'd230317442;
array2[5669]=30'd231362949;
array2[5670]=30'd229266819;
array2[5671]=30'd231362949;
array2[5672]=30'd229266819;
array2[5673]=30'd231364996;
array2[5674]=30'd230317442;
array2[5675]=30'd231362949;
array2[5676]=30'd230317442;
array2[5677]=30'd229266819;
array2[5678]=30'd228212100;
array2[5679]=30'd228212100;
array2[5680]=30'd228216193;
array2[5681]=30'd231362949;
array2[5682]=30'd230317442;
array2[5683]=30'd231364996;
array2[5684]=30'd179916222;
array2[5685]=30'd737318494;
array2[5686]=30'd790726247;
array2[5687]=30'd790726247;
array2[5688]=30'd790726247;
array2[5689]=30'd790726247;
array2[5690]=30'd790726247;
array2[5691]=30'd790726247;
array2[5692]=30'd764529268;
array2[5693]=30'd646130287;
array2[5694]=30'd646130287;
array2[5695]=30'd401997362;
array2[5696]=30'd179916222;
array2[5697]=30'd220861839;
array2[5698]=30'd227165569;
array2[5699]=30'd234504581;
array2[5700]=30'd231362949;
array2[5701]=30'd228216193;
array2[5702]=30'd227165569;
array2[5703]=30'd231364996;
array2[5704]=30'd229266819;
array2[5705]=30'd232417668;
array2[5706]=30'd225072515;
array2[5707]=30'd230317442;
array2[5708]=30'd230317442;
array2[5709]=30'd229266819;
array2[5710]=30'd229266819;
array2[5711]=30'd229266819;
array2[5712]=30'd229266819;
array2[5713]=30'd229266819;
array2[5714]=30'd231362949;
array2[5715]=30'd231364996;
array2[5716]=30'd231362949;
array2[5717]=30'd231359873;
array2[5718]=30'd231362949;
array2[5719]=30'd231364996;
array2[5720]=30'd230317442;
array2[5721]=30'd230317442;
array2[5722]=30'd229266819;
array2[5723]=30'd231362949;
array2[5724]=30'd231362949;
array2[5725]=30'd230317442;
array2[5726]=30'd231362949;
array2[5727]=30'd231362949;
array2[5728]=30'd230317442;
array2[5729]=30'd231362949;
array2[5730]=30'd230317442;
array2[5731]=30'd229266819;
array2[5732]=30'd231364996;
array2[5733]=30'd231362949;
array2[5734]=30'd229266819;
array2[5735]=30'd231362949;
array2[5736]=30'd229266819;
array2[5737]=30'd229266819;
array2[5738]=30'd230317442;
array2[5739]=30'd231362949;
array2[5740]=30'd228216193;
array2[5741]=30'd231362949;
array2[5742]=30'd230317442;
array2[5743]=30'd231362949;
array2[5744]=30'd231362949;
array2[5745]=30'd231364996;
array2[5746]=30'd231362949;
array2[5747]=30'd231362949;
array2[5748]=30'd231364996;
array2[5749]=30'd230317442;
array2[5750]=30'd234504581;
array2[5751]=30'd231364996;
array2[5752]=30'd231364996;
array2[5753]=30'd231364996;
array2[5754]=30'd231362949;
array2[5755]=30'd229266819;
array2[5756]=30'd229266819;
array2[5757]=30'd231362949;
array2[5758]=30'd229266819;
array2[5759]=30'd231362949;
array2[5760]=30'd193577377;
array2[5761]=30'd234504581;
array2[5762]=30'd227165569;
array2[5763]=30'd228216193;
array2[5764]=30'd230317442;
array2[5765]=30'd272255371;
array2[5766]=30'd401193372;
array2[5767]=30'd256519562;
array2[5768]=30'd229270912;
array2[5769]=30'd377085336;
array2[5770]=30'd603537847;
array2[5771]=30'd338288022;
array2[5772]=30'd231364996;
array2[5773]=30'd231364996;
array2[5774]=30'd231362949;
array2[5775]=30'd231364996;
array2[5776]=30'd230317442;
array2[5777]=30'd272255371;
array2[5778]=30'd553231776;
array2[5779]=30'd401193372;
array2[5780]=30'd179916222;
array2[5781]=30'd678604396;
array2[5782]=30'd764529268;
array2[5783]=30'd790726247;
array2[5784]=30'd790726247;
array2[5785]=30'd790726247;
array2[5786]=30'd790726247;
array2[5787]=30'd764529268;
array2[5788]=30'd790726247;
array2[5789]=30'd790726247;
array2[5790]=30'd790726247;
array2[5791]=30'd708987491;
array2[5792]=30'd646130287;
array2[5793]=30'd383147560;
array2[5794]=30'd260631016;
array2[5795]=30'd260631016;
array2[5796]=30'd220861839;
array2[5797]=30'd230307208;
array2[5798]=30'd228216193;
array2[5799]=30'd230317442;
array2[5800]=30'd227159434;
array2[5801]=30'd553231776;
array2[5802]=30'd472496545;
array2[5803]=30'd232392085;
array2[5804]=30'd231364996;
array2[5805]=30'd229266819;
array2[5806]=30'd231362949;
array2[5807]=30'd229266819;
array2[5808]=30'd231364996;
array2[5809]=30'd229266819;
array2[5810]=30'd231362949;
array2[5811]=30'd228216193;
array2[5812]=30'd231362949;
array2[5813]=30'd231362949;
array2[5814]=30'd231362949;
array2[5815]=30'd229266819;
array2[5816]=30'd229266819;
array2[5817]=30'd229266819;
array2[5818]=30'd229266819;
array2[5819]=30'd231362949;
array2[5820]=30'd231362949;
array2[5821]=30'd228216193;
array2[5822]=30'd231362949;
array2[5823]=30'd231362949;
array2[5824]=30'd231362949;
array2[5825]=30'd229266819;
array2[5826]=30'd231362949;
array2[5827]=30'd231362949;
array2[5828]=30'd231362949;
array2[5829]=30'd230317442;
array2[5830]=30'd231362949;
array2[5831]=30'd229266819;
array2[5832]=30'd231362949;
array2[5833]=30'd231362949;
array2[5834]=30'd229266819;
array2[5835]=30'd231362949;
array2[5836]=30'd229266819;
array2[5837]=30'd230317442;
array2[5838]=30'd231362949;
array2[5839]=30'd231362949;
array2[5840]=30'd231362949;
array2[5841]=30'd231362949;
array2[5842]=30'd231362949;
array2[5843]=30'd231362949;
array2[5844]=30'd231362949;
array2[5845]=30'd228216193;
array2[5846]=30'd231362949;
array2[5847]=30'd231362949;
array2[5848]=30'd230317442;
array2[5849]=30'd231364996;
array2[5850]=30'd229266819;
array2[5851]=30'd231362949;
array2[5852]=30'd230317442;
array2[5853]=30'd229266819;
array2[5854]=30'd231362949;
array2[5855]=30'd231364996;
array2[5856]=30'd193577377;
array2[5857]=30'd231359873;
array2[5858]=30'd227165569;
array2[5859]=30'd228216193;
array2[5860]=30'd230317442;
array2[5861]=30'd272255371;
array2[5862]=30'd377085336;
array2[5863]=30'd232422779;
array2[5864]=30'd231364996;
array2[5865]=30'd338288022;
array2[5866]=30'd532258209;
array2[5867]=30'd338288022;
array2[5868]=30'd229266819;
array2[5869]=30'd229266819;
array2[5870]=30'd231362949;
array2[5871]=30'd231362949;
array2[5872]=30'd231362949;
array2[5873]=30'd256519562;
array2[5874]=30'd472496545;
array2[5875]=30'd377085336;
array2[5876]=30'd179916222;
array2[5877]=30'd566515308;
array2[5878]=30'd762499681;
array2[5879]=30'd790726247;
array2[5880]=30'd790726247;
array2[5881]=30'd790726247;
array2[5882]=30'd790726247;
array2[5883]=30'd764529268;
array2[5884]=30'd790726247;
array2[5885]=30'd805398138;
array2[5886]=30'd790726247;
array2[5887]=30'd790726247;
array2[5888]=30'd764529268;
array2[5889]=30'd762499681;
array2[5890]=30'd727851632;
array2[5891]=30'd565444213;
array2[5892]=30'd249001484;
array2[5893]=30'd186252693;
array2[5894]=30'd229266819;
array2[5895]=30'd231364996;
array2[5896]=30'd231364996;
array2[5897]=30'd489282972;
array2[5898]=30'd464076202;
array2[5899]=30'd221916546;
array2[5900]=30'd227165569;
array2[5901]=30'd231362949;
array2[5902]=30'd229266819;
array2[5903]=30'd231362949;
array2[5904]=30'd231359873;
array2[5905]=30'd231362949;
array2[5906]=30'd231362949;
array2[5907]=30'd231362949;
array2[5908]=30'd228216193;
array2[5909]=30'd231362949;
array2[5910]=30'd231362949;
array2[5911]=30'd231359873;
array2[5912]=30'd229266819;
array2[5913]=30'd230317442;
array2[5914]=30'd231362949;
array2[5915]=30'd231362949;
array2[5916]=30'd228216193;
array2[5917]=30'd229266819;
array2[5918]=30'd231362949;
array2[5919]=30'd231362949;
array2[5920]=30'd228216193;
array2[5921]=30'd228216193;
array2[5922]=30'd231362949;
array2[5923]=30'd231362949;
array2[5924]=30'd234504581;
array2[5925]=30'd231362949;
array2[5926]=30'd228216193;
array2[5927]=30'd229266819;
array2[5928]=30'd228216193;
array2[5929]=30'd231362949;
array2[5930]=30'd231362949;
array2[5931]=30'd229266819;
array2[5932]=30'd230317442;
array2[5933]=30'd231362949;
array2[5934]=30'd231359873;
array2[5935]=30'd230317442;
array2[5936]=30'd231362949;
array2[5937]=30'd231362949;
array2[5938]=30'd231362949;
array2[5939]=30'd228216193;
array2[5940]=30'd228216193;
array2[5941]=30'd229266819;
array2[5942]=30'd229266819;
array2[5943]=30'd231362949;
array2[5944]=30'd228216193;
array2[5945]=30'd229266819;
array2[5946]=30'd231362949;
array2[5947]=30'd231362949;
array2[5948]=30'd228216193;
array2[5949]=30'd227165569;
array2[5950]=30'd228216193;
array2[5951]=30'd229266819;
array2[5952]=30'd193577377;
array2[5953]=30'd231359873;
array2[5954]=30'd227165569;
array2[5955]=30'd228216193;
array2[5956]=30'd230317442;
array2[5957]=30'd231362949;
array2[5958]=30'd229266819;
array2[5959]=30'd229270912;
array2[5960]=30'd232417668;
array2[5961]=30'd229266819;
array2[5962]=30'd228212100;
array2[5963]=30'd228216193;
array2[5964]=30'd231362949;
array2[5965]=30'd229266819;
array2[5966]=30'd231364996;
array2[5967]=30'd231364996;
array2[5968]=30'd229266819;
array2[5969]=30'd238691720;
array2[5970]=30'd227159434;
array2[5971]=30'd221916546;
array2[5972]=30'd240774546;
array2[5973]=30'd249001484;
array2[5974]=30'd737318494;
array2[5975]=30'd790726247;
array2[5976]=30'd790726247;
array2[5977]=30'd790726247;
array2[5978]=30'd790726247;
array2[5979]=30'd790726247;
array2[5980]=30'd790726247;
array2[5981]=30'd790726247;
array2[5982]=30'd790726247;
array2[5983]=30'd790726247;
array2[5984]=30'd790726247;
array2[5985]=30'd790726247;
array2[5986]=30'd790726247;
array2[5987]=30'd764529268;
array2[5988]=30'd483727963;
array2[5989]=30'd193577377;
array2[5990]=30'd228216193;
array2[5991]=30'd229266819;
array2[5992]=30'd231364996;
array2[5993]=30'd231364996;
array2[5994]=30'd227165569;
array2[5995]=30'd227165569;
array2[5996]=30'd229266819;
array2[5997]=30'd231362949;
array2[5998]=30'd231362949;
array2[5999]=30'd230317442;
array2[6000]=30'd228216193;
array2[6001]=30'd229266819;
array2[6002]=30'd229266819;
array2[6003]=30'd231362949;
array2[6004]=30'd234504581;
array2[6005]=30'd227165569;
array2[6006]=30'd229266819;
array2[6007]=30'd228216193;
array2[6008]=30'd231362949;
array2[6009]=30'd234504581;
array2[6010]=30'd231362949;
array2[6011]=30'd228216193;
array2[6012]=30'd228216193;
array2[6013]=30'd231362949;
array2[6014]=30'd231362949;
array2[6015]=30'd231362949;
array2[6016]=30'd231362949;
array2[6017]=30'd229266819;
array2[6018]=30'd229266819;
array2[6019]=30'd229266819;
array2[6020]=30'd231359873;
array2[6021]=30'd231364996;
array2[6022]=30'd231362949;
array2[6023]=30'd229266819;
array2[6024]=30'd228216193;
array2[6025]=30'd231362949;
array2[6026]=30'd231362949;
array2[6027]=30'd230317442;
array2[6028]=30'd229266819;
array2[6029]=30'd229266819;
array2[6030]=30'd231362949;
array2[6031]=30'd231362949;
array2[6032]=30'd229266819;
array2[6033]=30'd231362949;
array2[6034]=30'd231364996;
array2[6035]=30'd231362949;
array2[6036]=30'd229266819;
array2[6037]=30'd230317442;
array2[6038]=30'd231362949;
array2[6039]=30'd231362949;
array2[6040]=30'd229266819;
array2[6041]=30'd229266819;
array2[6042]=30'd231362949;
array2[6043]=30'd229266819;
array2[6044]=30'd231362949;
array2[6045]=30'd231362949;
array2[6046]=30'd227165569;
array2[6047]=30'd231364996;
array2[6048]=30'd193577377;
array2[6049]=30'd231359873;
array2[6050]=30'd227165569;
array2[6051]=30'd228216193;
array2[6052]=30'd230317442;
array2[6053]=30'd231362949;
array2[6054]=30'd229266819;
array2[6055]=30'd229270912;
array2[6056]=30'd234515845;
array2[6057]=30'd229266819;
array2[6058]=30'd231362949;
array2[6059]=30'd231362949;
array2[6060]=30'd229266819;
array2[6061]=30'd256519562;
array2[6062]=30'd532258209;
array2[6063]=30'd338288022;
array2[6064]=30'd225072515;
array2[6065]=30'd265928088;
array2[6066]=30'd280599950;
array2[6067]=30'd304706973;
array2[6068]=30'd304706973;
array2[6069]=30'd281508345;
array2[6070]=30'd727851632;
array2[6071]=30'd805398138;
array2[6072]=30'd823228019;
array2[6073]=30'd790726247;
array2[6074]=30'd805398138;
array2[6075]=30'd790726247;
array2[6076]=30'd790726247;
array2[6077]=30'd764529268;
array2[6078]=30'd790726247;
array2[6079]=30'd790726247;
array2[6080]=30'd790726247;
array2[6081]=30'd790726247;
array2[6082]=30'd790726247;
array2[6083]=30'd727851632;
array2[6084]=30'd407216718;
array2[6085]=30'd464076202;
array2[6086]=30'd425297329;
array2[6087]=30'd234515845;
array2[6088]=30'd229266819;
array2[6089]=30'd236604812;
array2[6090]=30'd227165569;
array2[6091]=30'd229266819;
array2[6092]=30'd231364996;
array2[6093]=30'd231362949;
array2[6094]=30'd231362949;
array2[6095]=30'd230317442;
array2[6096]=30'd231364996;
array2[6097]=30'd231362949;
array2[6098]=30'd231362949;
array2[6099]=30'd229266819;
array2[6100]=30'd228216193;
array2[6101]=30'd231362949;
array2[6102]=30'd229266819;
array2[6103]=30'd231359873;
array2[6104]=30'd231359873;
array2[6105]=30'd227165569;
array2[6106]=30'd229266819;
array2[6107]=30'd234504581;
array2[6108]=30'd234504581;
array2[6109]=30'd228216193;
array2[6110]=30'd229266819;
array2[6111]=30'd231362949;
array2[6112]=30'd234504581;
array2[6113]=30'd231362949;
array2[6114]=30'd229266819;
array2[6115]=30'd229266819;
array2[6116]=30'd231362949;
array2[6117]=30'd229266819;
array2[6118]=30'd229266819;
array2[6119]=30'd229266819;
array2[6120]=30'd229266819;
array2[6121]=30'd231362949;
array2[6122]=30'd229266819;
array2[6123]=30'd231362949;
array2[6124]=30'd231362949;
array2[6125]=30'd231362949;
array2[6126]=30'd231362949;
array2[6127]=30'd230317442;
array2[6128]=30'd229266819;
array2[6129]=30'd229266819;
array2[6130]=30'd231362949;
array2[6131]=30'd229266819;
array2[6132]=30'd229266819;
array2[6133]=30'd234504581;
array2[6134]=30'd231364996;
array2[6135]=30'd231362949;
array2[6136]=30'd231362949;
array2[6137]=30'd229266819;
array2[6138]=30'd231362949;
array2[6139]=30'd231362949;
array2[6140]=30'd231362949;
array2[6141]=30'd231362949;
array2[6142]=30'd229266819;
array2[6143]=30'd229266819;
array2[6144]=30'd193577377;
array2[6145]=30'd231359873;
array2[6146]=30'd227165569;
array2[6147]=30'd228216193;
array2[6148]=30'd230317442;
array2[6149]=30'd231362949;
array2[6150]=30'd229266819;
array2[6151]=30'd229270912;
array2[6152]=30'd234515845;
array2[6153]=30'd229266819;
array2[6154]=30'd231362949;
array2[6155]=30'd231362949;
array2[6156]=30'd231362949;
array2[6157]=30'd272255371;
array2[6158]=30'd553231776;
array2[6159]=30'd338288022;
array2[6160]=30'd230317442;
array2[6161]=30'd262793620;
array2[6162]=30'd280599950;
array2[6163]=30'd312021416;
array2[6164]=30'd280599950;
array2[6165]=30'd281508345;
array2[6166]=30'd450208341;
array2[6167]=30'd483727963;
array2[6168]=30'd506770009;
array2[6169]=30'd483727963;
array2[6170]=30'd678602388;
array2[6171]=30'd764529268;
array2[6172]=30'd805398138;
array2[6173]=30'd790726247;
array2[6174]=30'd790726247;
array2[6175]=30'd790726247;
array2[6176]=30'd790726247;
array2[6177]=30'd790726247;
array2[6178]=30'd790726247;
array2[6179]=30'd645112409;
array2[6180]=30'd207191473;
array2[6181]=30'd532258209;
array2[6182]=30'd405404052;
array2[6183]=30'd231362949;
array2[6184]=30'd229266819;
array2[6185]=30'd232417668;
array2[6186]=30'd227165569;
array2[6187]=30'd230317442;
array2[6188]=30'd231362949;
array2[6189]=30'd231362949;
array2[6190]=30'd229266819;
array2[6191]=30'd229266819;
array2[6192]=30'd231362949;
array2[6193]=30'd231359873;
array2[6194]=30'd231362949;
array2[6195]=30'd231362949;
array2[6196]=30'd230317442;
array2[6197]=30'd231362949;
array2[6198]=30'd231359873;
array2[6199]=30'd229266819;
array2[6200]=30'd231362949;
array2[6201]=30'd229266819;
array2[6202]=30'd230317442;
array2[6203]=30'd231362949;
array2[6204]=30'd231362949;
array2[6205]=30'd231359873;
array2[6206]=30'd229266819;
array2[6207]=30'd228216193;
array2[6208]=30'd234504581;
array2[6209]=30'd231362949;
array2[6210]=30'd228216193;
array2[6211]=30'd229266819;
array2[6212]=30'd228216193;
array2[6213]=30'd231362949;
array2[6214]=30'd234504581;
array2[6215]=30'd227165569;
array2[6216]=30'd231362949;
array2[6217]=30'd231362949;
array2[6218]=30'd231364996;
array2[6219]=30'd231362949;
array2[6220]=30'd231362949;
array2[6221]=30'd230317442;
array2[6222]=30'd231362949;
array2[6223]=30'd231364996;
array2[6224]=30'd231364996;
array2[6225]=30'd229266819;
array2[6226]=30'd228216193;
array2[6227]=30'd231362949;
array2[6228]=30'd229266819;
array2[6229]=30'd234504581;
array2[6230]=30'd228216193;
array2[6231]=30'd228216193;
array2[6232]=30'd231359873;
array2[6233]=30'd231362949;
array2[6234]=30'd231362949;
array2[6235]=30'd231362949;
array2[6236]=30'd229266819;
array2[6237]=30'd231362949;
array2[6238]=30'd231362949;
array2[6239]=30'd229266819;
array2[6240]=30'd193577377;
array2[6241]=30'd234504581;
array2[6242]=30'd227165569;
array2[6243]=30'd228216193;
array2[6244]=30'd230317442;
array2[6245]=30'd231362949;
array2[6246]=30'd229266819;
array2[6247]=30'd229270912;
array2[6248]=30'd234515845;
array2[6249]=30'd229266819;
array2[6250]=30'd231362949;
array2[6251]=30'd229270912;
array2[6252]=30'd231362949;
array2[6253]=30'd231362949;
array2[6254]=30'd229266819;
array2[6255]=30'd230317442;
array2[6256]=30'd231364996;
array2[6257]=30'd240774546;
array2[6258]=30'd304706973;
array2[6259]=30'd295249323;
array2[6260]=30'd304706973;
array2[6261]=30'd254365107;
array2[6262]=30'd254365107;
array2[6263]=30'd254365107;
array2[6264]=30'd254365107;
array2[6265]=30'd254365107;
array2[6266]=30'd383147560;
array2[6267]=30'd407216718;
array2[6268]=30'd444954173;
array2[6269]=30'd407216718;
array2[6270]=30'd566515308;
array2[6271]=30'd764529268;
array2[6272]=30'd790726247;
array2[6273]=30'd790726247;
array2[6274]=30'd708987491;
array2[6275]=30'd319215128;
array2[6276]=30'd212454818;
array2[6277]=30'd227165569;
array2[6278]=30'd231362949;
array2[6279]=30'd228212100;
array2[6280]=30'd231362949;
array2[6281]=30'd231362949;
array2[6282]=30'd231362949;
array2[6283]=30'd229270912;
array2[6284]=30'd228216193;
array2[6285]=30'd230317442;
array2[6286]=30'd228216193;
array2[6287]=30'd231362949;
array2[6288]=30'd231362949;
array2[6289]=30'd231362949;
array2[6290]=30'd230317442;
array2[6291]=30'd231362949;
array2[6292]=30'd230317442;
array2[6293]=30'd231362949;
array2[6294]=30'd230317442;
array2[6295]=30'd231362949;
array2[6296]=30'd230317442;
array2[6297]=30'd229266819;
array2[6298]=30'd230317442;
array2[6299]=30'd229266819;
array2[6300]=30'd229266819;
array2[6301]=30'd231362949;
array2[6302]=30'd229266819;
array2[6303]=30'd231362949;
array2[6304]=30'd231364996;
array2[6305]=30'd231362949;
array2[6306]=30'd230317442;
array2[6307]=30'd231362949;
array2[6308]=30'd229266819;
array2[6309]=30'd231362949;
array2[6310]=30'd231362949;
array2[6311]=30'd230317442;
array2[6312]=30'd234504581;
array2[6313]=30'd231364996;
array2[6314]=30'd231362949;
array2[6315]=30'd231362949;
array2[6316]=30'd230317442;
array2[6317]=30'd229266819;
array2[6318]=30'd228216193;
array2[6319]=30'd231359873;
array2[6320]=30'd231362949;
array2[6321]=30'd231362949;
array2[6322]=30'd229266819;
array2[6323]=30'd228216193;
array2[6324]=30'd231362949;
array2[6325]=30'd231359873;
array2[6326]=30'd231362949;
array2[6327]=30'd231362949;
array2[6328]=30'd231362949;
array2[6329]=30'd229266819;
array2[6330]=30'd231362949;
array2[6331]=30'd231362949;
array2[6332]=30'd231362949;
array2[6333]=30'd229266819;
array2[6334]=30'd228216193;
array2[6335]=30'd231362949;
array2[6336]=30'd193577377;
array2[6337]=30'd231359873;
array2[6338]=30'd227165569;
array2[6339]=30'd228216193;
array2[6340]=30'd230317442;
array2[6341]=30'd231362949;
array2[6342]=30'd229266819;
array2[6343]=30'd229270912;
array2[6344]=30'd234515845;
array2[6345]=30'd229266819;
array2[6346]=30'd231362949;
array2[6347]=30'd234515845;
array2[6348]=30'd231362949;
array2[6349]=30'd229266819;
array2[6350]=30'd229270912;
array2[6351]=30'd227165569;
array2[6352]=30'd231362949;
array2[6353]=30'd238691720;
array2[6354]=30'd304706973;
array2[6355]=30'd295249323;
array2[6356]=30'd312021416;
array2[6357]=30'd312021416;
array2[6358]=30'd304706973;
array2[6359]=30'd312021416;
array2[6360]=30'd312021416;
array2[6361]=30'd312021416;
array2[6362]=30'd312021416;
array2[6363]=30'd312021416;
array2[6364]=30'd312021416;
array2[6365]=30'd295249323;
array2[6366]=30'd260631016;
array2[6367]=30'd645112409;
array2[6368]=30'd790726247;
array2[6369]=30'd790726247;
array2[6370]=30'd678604396;
array2[6371]=30'd179916222;
array2[6372]=30'd227165569;
array2[6373]=30'd229266819;
array2[6374]=30'd229266819;
array2[6375]=30'd231362949;
array2[6376]=30'd231362949;
array2[6377]=30'd231362949;
array2[6378]=30'd231362949;
array2[6379]=30'd231364996;
array2[6380]=30'd229266819;
array2[6381]=30'd231362949;
array2[6382]=30'd229266819;
array2[6383]=30'd229266819;
array2[6384]=30'd231362949;
array2[6385]=30'd229266819;
array2[6386]=30'd229266819;
array2[6387]=30'd231362949;
array2[6388]=30'd231362949;
array2[6389]=30'd230317442;
array2[6390]=30'd230317442;
array2[6391]=30'd231362949;
array2[6392]=30'd231362949;
array2[6393]=30'd231364996;
array2[6394]=30'd230317442;
array2[6395]=30'd231362949;
array2[6396]=30'd231362949;
array2[6397]=30'd231362949;
array2[6398]=30'd231362949;
array2[6399]=30'd229266819;
array2[6400]=30'd231364996;
array2[6401]=30'd229266819;
array2[6402]=30'd229266819;
array2[6403]=30'd231362949;
array2[6404]=30'd231364996;
array2[6405]=30'd231362949;
array2[6406]=30'd230317442;
array2[6407]=30'd231362949;
array2[6408]=30'd229266819;
array2[6409]=30'd231362949;
array2[6410]=30'd230317442;
array2[6411]=30'd229266819;
array2[6412]=30'd231362949;
array2[6413]=30'd231364996;
array2[6414]=30'd231362949;
array2[6415]=30'd231362949;
array2[6416]=30'd229266819;
array2[6417]=30'd231362949;
array2[6418]=30'd229266819;
array2[6419]=30'd229266819;
array2[6420]=30'd228216193;
array2[6421]=30'd228216193;
array2[6422]=30'd230317442;
array2[6423]=30'd231362949;
array2[6424]=30'd231362949;
array2[6425]=30'd231364996;
array2[6426]=30'd231359873;
array2[6427]=30'd231362949;
array2[6428]=30'd230317442;
array2[6429]=30'd229266819;
array2[6430]=30'd231362949;
array2[6431]=30'd227165569;
array2[6432]=30'd193577377;
array2[6433]=30'd234504581;
array2[6434]=30'd227165569;
array2[6435]=30'd228216193;
array2[6436]=30'd230317442;
array2[6437]=30'd231362949;
array2[6438]=30'd229266819;
array2[6439]=30'd229270912;
array2[6440]=30'd234515845;
array2[6441]=30'd229266819;
array2[6442]=30'd231362949;
array2[6443]=30'd234515845;
array2[6444]=30'd230317442;
array2[6445]=30'd231362949;
array2[6446]=30'd231362949;
array2[6447]=30'd231364996;
array2[6448]=30'd230317442;
array2[6449]=30'd238691720;
array2[6450]=30'd304706973;
array2[6451]=30'd312021416;
array2[6452]=30'd312021416;
array2[6453]=30'd312021416;
array2[6454]=30'd304706973;
array2[6455]=30'd304706973;
array2[6456]=30'd312021416;
array2[6457]=30'd295249323;
array2[6458]=30'd304706973;
array2[6459]=30'd312021416;
array2[6460]=30'd304706973;
array2[6461]=30'd312021416;
array2[6462]=30'd195647926;
array2[6463]=30'd645112409;
array2[6464]=30'd790726247;
array2[6465]=30'd764529268;
array2[6466]=30'd565444213;
array2[6467]=30'd179916222;
array2[6468]=30'd231362949;
array2[6469]=30'd234504581;
array2[6470]=30'd231362949;
array2[6471]=30'd231362949;
array2[6472]=30'd230317442;
array2[6473]=30'd231362949;
array2[6474]=30'd230317442;
array2[6475]=30'd231362949;
array2[6476]=30'd230317442;
array2[6477]=30'd229266819;
array2[6478]=30'd229266819;
array2[6479]=30'd231362949;
array2[6480]=30'd229266819;
array2[6481]=30'd231362949;
array2[6482]=30'd231362949;
array2[6483]=30'd231362949;
array2[6484]=30'd231364996;
array2[6485]=30'd231362949;
array2[6486]=30'd230317442;
array2[6487]=30'd229266819;
array2[6488]=30'd231362949;
array2[6489]=30'd229266819;
array2[6490]=30'd231362949;
array2[6491]=30'd231362949;
array2[6492]=30'd231362949;
array2[6493]=30'd231362949;
array2[6494]=30'd231364996;
array2[6495]=30'd231362949;
array2[6496]=30'd230317442;
array2[6497]=30'd231362949;
array2[6498]=30'd231362949;
array2[6499]=30'd228216193;
array2[6500]=30'd230317442;
array2[6501]=30'd231364996;
array2[6502]=30'd231362949;
array2[6503]=30'd229266819;
array2[6504]=30'd230317442;
array2[6505]=30'd231362949;
array2[6506]=30'd231362949;
array2[6507]=30'd229266819;
array2[6508]=30'd229266819;
array2[6509]=30'd228216193;
array2[6510]=30'd231362949;
array2[6511]=30'd231362949;
array2[6512]=30'd231359873;
array2[6513]=30'd227165569;
array2[6514]=30'd231362949;
array2[6515]=30'd231362949;
array2[6516]=30'd231364996;
array2[6517]=30'd228216193;
array2[6518]=30'd229266819;
array2[6519]=30'd231362949;
array2[6520]=30'd231362949;
array2[6521]=30'd231362949;
array2[6522]=30'd234504581;
array2[6523]=30'd231364996;
array2[6524]=30'd231364996;
array2[6525]=30'd230317442;
array2[6526]=30'd231362949;
array2[6527]=30'd229266819;
array2[6528]=30'd193577377;
array2[6529]=30'd234504581;
array2[6530]=30'd227165569;
array2[6531]=30'd228216193;
array2[6532]=30'd229266819;
array2[6533]=30'd229266819;
array2[6534]=30'd229266819;
array2[6535]=30'd230317442;
array2[6536]=30'd230317442;
array2[6537]=30'd229266819;
array2[6538]=30'd231362949;
array2[6539]=30'd232417668;
array2[6540]=30'd231362949;
array2[6541]=30'd231362949;
array2[6542]=30'd229266819;
array2[6543]=30'd231364996;
array2[6544]=30'd230317442;
array2[6545]=30'd221916546;
array2[6546]=30'd304706973;
array2[6547]=30'd295249323;
array2[6548]=30'd312021416;
array2[6549]=30'd312021416;
array2[6550]=30'd312021416;
array2[6551]=30'd312021416;
array2[6552]=30'd312021416;
array2[6553]=30'd304706973;
array2[6554]=30'd295249323;
array2[6555]=30'd304706973;
array2[6556]=30'd312021416;
array2[6557]=30'd295249323;
array2[6558]=30'd195647926;
array2[6559]=30'd645112409;
array2[6560]=30'd790726247;
array2[6561]=30'd729975381;
array2[6562]=30'd190356956;
array2[6563]=30'd193577377;
array2[6564]=30'd212454818;
array2[6565]=30'd213516691;
array2[6566]=30'd236604812;
array2[6567]=30'd228216193;
array2[6568]=30'd231362949;
array2[6569]=30'd230317442;
array2[6570]=30'd231359873;
array2[6571]=30'd229266819;
array2[6572]=30'd231362949;
array2[6573]=30'd231362949;
array2[6574]=30'd231362949;
array2[6575]=30'd231362949;
array2[6576]=30'd229266819;
array2[6577]=30'd231362949;
array2[6578]=30'd230317442;
array2[6579]=30'd229266819;
array2[6580]=30'd231362949;
array2[6581]=30'd229266819;
array2[6582]=30'd231362949;
array2[6583]=30'd231362949;
array2[6584]=30'd231362949;
array2[6585]=30'd231362949;
array2[6586]=30'd228216193;
array2[6587]=30'd234504581;
array2[6588]=30'd231364996;
array2[6589]=30'd231362949;
array2[6590]=30'd229266819;
array2[6591]=30'd227165569;
array2[6592]=30'd231362949;
array2[6593]=30'd231362949;
array2[6594]=30'd234504581;
array2[6595]=30'd231364996;
array2[6596]=30'd231362949;
array2[6597]=30'd231362949;
array2[6598]=30'd231364996;
array2[6599]=30'd229266819;
array2[6600]=30'd229266819;
array2[6601]=30'd231362949;
array2[6602]=30'd229266819;
array2[6603]=30'd229266819;
array2[6604]=30'd230317442;
array2[6605]=30'd229266819;
array2[6606]=30'd231364996;
array2[6607]=30'd231362949;
array2[6608]=30'd229266819;
array2[6609]=30'd231362949;
array2[6610]=30'd230317442;
array2[6611]=30'd231362949;
array2[6612]=30'd230317442;
array2[6613]=30'd231362949;
array2[6614]=30'd229266819;
array2[6615]=30'd231362949;
array2[6616]=30'd231362949;
array2[6617]=30'd231362949;
array2[6618]=30'd231362949;
array2[6619]=30'd231364996;
array2[6620]=30'd231362949;
array2[6621]=30'd229266819;
array2[6622]=30'd231364996;
array2[6623]=30'd229266819;
array2[6624]=30'd193577377;
array2[6625]=30'd234504581;
array2[6626]=30'd227165569;
array2[6627]=30'd228216193;
array2[6628]=30'd230317442;
array2[6629]=30'd230317442;
array2[6630]=30'd229266819;
array2[6631]=30'd229270912;
array2[6632]=30'd229270912;
array2[6633]=30'd229266819;
array2[6634]=30'd231362949;
array2[6635]=30'd232417668;
array2[6636]=30'd229266819;
array2[6637]=30'd231362949;
array2[6638]=30'd229266819;
array2[6639]=30'd230317442;
array2[6640]=30'd231362949;
array2[6641]=30'd234504581;
array2[6642]=30'd262793620;
array2[6643]=30'd262793620;
array2[6644]=30'd265928088;
array2[6645]=30'd269069720;
array2[6646]=30'd265928088;
array2[6647]=30'd265928088;
array2[6648]=30'd280599950;
array2[6649]=30'd312021416;
array2[6650]=30'd312021416;
array2[6651]=30'd304706973;
array2[6652]=30'd312021416;
array2[6653]=30'd295249323;
array2[6654]=30'd190356956;
array2[6655]=30'd645112409;
array2[6656]=30'd790726247;
array2[6657]=30'd749877860;
array2[6658]=30'd483727963;
array2[6659]=30'd450208341;
array2[6660]=30'd319215128;
array2[6661]=30'd179916222;
array2[6662]=30'd193577377;
array2[6663]=30'd232392085;
array2[6664]=30'd231364996;
array2[6665]=30'd231362949;
array2[6666]=30'd230317442;
array2[6667]=30'd229266819;
array2[6668]=30'd231362949;
array2[6669]=30'd229266819;
array2[6670]=30'd231362949;
array2[6671]=30'd231362949;
array2[6672]=30'd231362949;
array2[6673]=30'd229266819;
array2[6674]=30'd236604812;
array2[6675]=30'd256519562;
array2[6676]=30'd256519562;
array2[6677]=30'd229266819;
array2[6678]=30'd229266819;
array2[6679]=30'd229266819;
array2[6680]=30'd231362949;
array2[6681]=30'd231362949;
array2[6682]=30'd234504581;
array2[6683]=30'd229266819;
array2[6684]=30'd231362949;
array2[6685]=30'd231362949;
array2[6686]=30'd231362949;
array2[6687]=30'd272255371;
array2[6688]=30'd338288022;
array2[6689]=30'd231364996;
array2[6690]=30'd228216193;
array2[6691]=30'd229266819;
array2[6692]=30'd228216193;
array2[6693]=30'd231364996;
array2[6694]=30'd231362949;
array2[6695]=30'd229266819;
array2[6696]=30'd231362949;
array2[6697]=30'd230317442;
array2[6698]=30'd231362949;
array2[6699]=30'd230317442;
array2[6700]=30'd229266819;
array2[6701]=30'd230317442;
array2[6702]=30'd231362949;
array2[6703]=30'd229266819;
array2[6704]=30'd229266819;
array2[6705]=30'd231362949;
array2[6706]=30'd231362949;
array2[6707]=30'd230317442;
array2[6708]=30'd231362949;
array2[6709]=30'd229266819;
array2[6710]=30'd231362949;
array2[6711]=30'd231364996;
array2[6712]=30'd231362949;
array2[6713]=30'd231364996;
array2[6714]=30'd231362949;
array2[6715]=30'd231362949;
array2[6716]=30'd231362949;
array2[6717]=30'd230317442;
array2[6718]=30'd230317442;
array2[6719]=30'd231362949;
array2[6720]=30'd193577377;
array2[6721]=30'd234504581;
array2[6722]=30'd227165569;
array2[6723]=30'd228216193;
array2[6724]=30'd230317442;
array2[6725]=30'd231362949;
array2[6726]=30'd229266819;
array2[6727]=30'd229270912;
array2[6728]=30'd234515845;
array2[6729]=30'd229266819;
array2[6730]=30'd231362949;
array2[6731]=30'd234515845;
array2[6732]=30'd230317442;
array2[6733]=30'd231362949;
array2[6734]=30'd229266819;
array2[6735]=30'd231362949;
array2[6736]=30'd229266819;
array2[6737]=30'd231364996;
array2[6738]=30'd230317442;
array2[6739]=30'd229266819;
array2[6740]=30'd231362949;
array2[6741]=30'd227165569;
array2[6742]=30'd230307208;
array2[6743]=30'd234504581;
array2[6744]=30'd265928088;
array2[6745]=30'd265928088;
array2[6746]=30'd265928088;
array2[6747]=30'd265928088;
array2[6748]=30'd280599950;
array2[6749]=30'd254365107;
array2[6750]=30'd347490866;
array2[6751]=30'd678604396;
array2[6752]=30'd790726247;
array2[6753]=30'd790726247;
array2[6754]=30'd790726247;
array2[6755]=30'd764529268;
array2[6756]=30'd645112409;
array2[6757]=30'd506770009;
array2[6758]=30'd249001484;
array2[6759]=30'd220861839;
array2[6760]=30'd231364996;
array2[6761]=30'd231362949;
array2[6762]=30'd231362949;
array2[6763]=30'd231362949;
array2[6764]=30'd231362949;
array2[6765]=30'd231359873;
array2[6766]=30'd231362949;
array2[6767]=30'd231362949;
array2[6768]=30'd256519562;
array2[6769]=30'd236604812;
array2[6770]=30'd272255371;
array2[6771]=30'd428475791;
array2[6772]=30'd272255371;
array2[6773]=30'd234504581;
array2[6774]=30'd272255371;
array2[6775]=30'd228216193;
array2[6776]=30'd230307208;
array2[6777]=30'd227165569;
array2[6778]=30'd227165569;
array2[6779]=30'd227165569;
array2[6780]=30'd232392085;
array2[6781]=30'd227159434;
array2[6782]=30'd221916546;
array2[6783]=30'd603537847;
array2[6784]=30'd655981997;
array2[6785]=30'd256519562;
array2[6786]=30'd228216193;
array2[6787]=30'd231359873;
array2[6788]=30'd229266819;
array2[6789]=30'd229270912;
array2[6790]=30'd231364996;
array2[6791]=30'd228216193;
array2[6792]=30'd231359873;
array2[6793]=30'd229266819;
array2[6794]=30'd231362949;
array2[6795]=30'd231362949;
array2[6796]=30'd231362949;
array2[6797]=30'd231362949;
array2[6798]=30'd229266819;
array2[6799]=30'd231364996;
array2[6800]=30'd231364996;
array2[6801]=30'd229266819;
array2[6802]=30'd228216193;
array2[6803]=30'd229266819;
array2[6804]=30'd229266819;
array2[6805]=30'd231362949;
array2[6806]=30'd231362949;
array2[6807]=30'd231362949;
array2[6808]=30'd231362949;
array2[6809]=30'd231362949;
array2[6810]=30'd229266819;
array2[6811]=30'd231364996;
array2[6812]=30'd231364996;
array2[6813]=30'd231364996;
array2[6814]=30'd234504581;
array2[6815]=30'd229266819;
array2[6816]=30'd193577377;
array2[6817]=30'd231359873;
array2[6818]=30'd227165569;
array2[6819]=30'd228216193;
array2[6820]=30'd230317442;
array2[6821]=30'd231362949;
array2[6822]=30'd229266819;
array2[6823]=30'd229270912;
array2[6824]=30'd234515845;
array2[6825]=30'd229266819;
array2[6826]=30'd231362949;
array2[6827]=30'd234515845;
array2[6828]=30'd230317442;
array2[6829]=30'd231362949;
array2[6830]=30'd229266819;
array2[6831]=30'd231359873;
array2[6832]=30'd229266819;
array2[6833]=30'd229266819;
array2[6834]=30'd231362949;
array2[6835]=30'd228216193;
array2[6836]=30'd231359873;
array2[6837]=30'd229266819;
array2[6838]=30'd231362949;
array2[6839]=30'd231362949;
array2[6840]=30'd234504581;
array2[6841]=30'd231362949;
array2[6842]=30'd231362949;
array2[6843]=30'd231362949;
array2[6844]=30'd271165847;
array2[6845]=30'd254365107;
array2[6846]=30'd265736724;
array2[6847]=30'd560184961;
array2[6848]=30'd762499681;
array2[6849]=30'd764529268;
array2[6850]=30'd764529268;
array2[6851]=30'd764529268;
array2[6852]=30'd764529268;
array2[6853]=30'd764529268;
array2[6854]=30'd319215128;
array2[6855]=30'd221916546;
array2[6856]=30'd231364996;
array2[6857]=30'd227165569;
array2[6858]=30'd229266819;
array2[6859]=30'd230317442;
array2[6860]=30'd230317442;
array2[6861]=30'd231362949;
array2[6862]=30'd229266819;
array2[6863]=30'd229266819;
array2[6864]=30'd401193372;
array2[6865]=30'd301610387;
array2[6866]=30'd229266819;
array2[6867]=30'd229270912;
array2[6868]=30'd228216193;
array2[6869]=30'd272255371;
array2[6870]=30'd401193372;
array2[6871]=30'd207191473;
array2[6872]=30'd150539724;
array2[6873]=30'd179916222;
array2[6874]=30'd232392085;
array2[6875]=30'd232392085;
array2[6876]=30'd257539480;
array2[6877]=30'd269069720;
array2[6878]=30'd228181405;
array2[6879]=30'd532258209;
array2[6880]=30'd532258209;
array2[6881]=30'd238691720;
array2[6882]=30'd231362949;
array2[6883]=30'd229266819;
array2[6884]=30'd231362949;
array2[6885]=30'd231364996;
array2[6886]=30'd230317442;
array2[6887]=30'd229266819;
array2[6888]=30'd231362949;
array2[6889]=30'd229266819;
array2[6890]=30'd229266819;
array2[6891]=30'd229266819;
array2[6892]=30'd231362949;
array2[6893]=30'd231362949;
array2[6894]=30'd229266819;
array2[6895]=30'd228216193;
array2[6896]=30'd228216193;
array2[6897]=30'd228216193;
array2[6898]=30'd228216193;
array2[6899]=30'd230317442;
array2[6900]=30'd230317442;
array2[6901]=30'd230317442;
array2[6902]=30'd231362949;
array2[6903]=30'd229266819;
array2[6904]=30'd230317442;
array2[6905]=30'd231362949;
array2[6906]=30'd231362949;
array2[6907]=30'd231362949;
array2[6908]=30'd231362949;
array2[6909]=30'd229266819;
array2[6910]=30'd227165569;
array2[6911]=30'd228216193;
array2[6912]=30'd193577377;
array2[6913]=30'd234504581;
array2[6914]=30'd227165569;
array2[6915]=30'd228216193;
array2[6916]=30'd230317442;
array2[6917]=30'd229266819;
array2[6918]=30'd229266819;
array2[6919]=30'd230317442;
array2[6920]=30'd229270912;
array2[6921]=30'd229266819;
array2[6922]=30'd231362949;
array2[6923]=30'd229270912;
array2[6924]=30'd230317442;
array2[6925]=30'd231362949;
array2[6926]=30'd229266819;
array2[6927]=30'd231359873;
array2[6928]=30'd229266819;
array2[6929]=30'd228216193;
array2[6930]=30'd229266819;
array2[6931]=30'd231362949;
array2[6932]=30'd231362949;
array2[6933]=30'd231362949;
array2[6934]=30'd231364996;
array2[6935]=30'd256519562;
array2[6936]=30'd256519562;
array2[6937]=30'd234504581;
array2[6938]=30'd231362949;
array2[6939]=30'd231362949;
array2[6940]=30'd304706973;
array2[6941]=30'd271165847;
array2[6942]=30'd207191473;
array2[6943]=30'd281508345;
array2[6944]=30'd319215128;
array2[6945]=30'd319215128;
array2[6946]=30'd319215128;
array2[6947]=30'd319215128;
array2[6948]=30'd566515308;
array2[6949]=30'd678604396;
array2[6950]=30'd281508345;
array2[6951]=30'd220861839;
array2[6952]=30'd231362949;
array2[6953]=30'd231364996;
array2[6954]=30'd231362949;
array2[6955]=30'd230317442;
array2[6956]=30'd231364996;
array2[6957]=30'd231362949;
array2[6958]=30'd229270912;
array2[6959]=30'd272255371;
array2[6960]=30'd236604812;
array2[6961]=30'd231362949;
array2[6962]=30'd231362949;
array2[6963]=30'd227165569;
array2[6964]=30'd213516691;
array2[6965]=30'd213516691;
array2[6966]=30'd234499470;
array2[6967]=30'd254365107;
array2[6968]=30'd124307934;
array2[6969]=30'd159912438;
array2[6970]=30'd190356956;
array2[6971]=30'd281508345;
array2[6972]=30'd260631016;
array2[6973]=30'd248105365;
array2[6974]=30'd269069720;
array2[6975]=30'd248105365;
array2[6976]=30'd240774546;
array2[6977]=30'd248105365;
array2[6978]=30'd238691720;
array2[6979]=30'd227165569;
array2[6980]=30'd227165569;
array2[6981]=30'd227165569;
array2[6982]=30'd231359873;
array2[6983]=30'd229266819;
array2[6984]=30'd231362949;
array2[6985]=30'd231362949;
array2[6986]=30'd231362949;
array2[6987]=30'd231362949;
array2[6988]=30'd231362949;
array2[6989]=30'd231362949;
array2[6990]=30'd231362949;
array2[6991]=30'd231362949;
array2[6992]=30'd231362949;
array2[6993]=30'd230317442;
array2[6994]=30'd229266819;
array2[6995]=30'd230317442;
array2[6996]=30'd231362949;
array2[6997]=30'd231362949;
array2[6998]=30'd231362949;
array2[6999]=30'd229266819;
array2[7000]=30'd229266819;
array2[7001]=30'd229266819;
array2[7002]=30'd229266819;
array2[7003]=30'd231362949;
array2[7004]=30'd231362949;
array2[7005]=30'd231362949;
array2[7006]=30'd229266819;
array2[7007]=30'd231362949;
array2[7008]=30'd193577377;
array2[7009]=30'd231359873;
array2[7010]=30'd227165569;
array2[7011]=30'd228216193;
array2[7012]=30'd230317442;
array2[7013]=30'd231362949;
array2[7014]=30'd229266819;
array2[7015]=30'd229270912;
array2[7016]=30'd234515845;
array2[7017]=30'd229266819;
array2[7018]=30'd231362949;
array2[7019]=30'd234515845;
array2[7020]=30'd230317442;
array2[7021]=30'd231362949;
array2[7022]=30'd229266819;
array2[7023]=30'd231359873;
array2[7024]=30'd229266819;
array2[7025]=30'd229266819;
array2[7026]=30'd229266819;
array2[7027]=30'd231362949;
array2[7028]=30'd231362949;
array2[7029]=30'd231362949;
array2[7030]=30'd231362949;
array2[7031]=30'd338288022;
array2[7032]=30'd301610387;
array2[7033]=30'd231362949;
array2[7034]=30'd234504581;
array2[7035]=30'd234504581;
array2[7036]=30'd304706973;
array2[7037]=30'd271165847;
array2[7038]=30'd221916546;
array2[7039]=30'd221916546;
array2[7040]=30'd232392085;
array2[7041]=30'd232392085;
array2[7042]=30'd227159434;
array2[7043]=30'd207191473;
array2[7044]=30'd299264555;
array2[7045]=30'd265736724;
array2[7046]=30'd228181405;
array2[7047]=30'd228212100;
array2[7048]=30'd228216193;
array2[7049]=30'd228216193;
array2[7050]=30'd231362949;
array2[7051]=30'd230317442;
array2[7052]=30'd230317442;
array2[7053]=30'd231362949;
array2[7054]=30'd301610387;
array2[7055]=30'd428475791;
array2[7056]=30'd256519562;
array2[7057]=30'd234504581;
array2[7058]=30'd228216193;
array2[7059]=30'd212454818;
array2[7060]=30'd124307934;
array2[7061]=30'd124307934;
array2[7062]=30'd179916222;
array2[7063]=30'd338288022;
array2[7064]=30'd190356956;
array2[7065]=30'd208120309;
array2[7066]=30'd347490866;
array2[7067]=30'd560184961;
array2[7068]=30'd449120871;
array2[7069]=30'd299264555;
array2[7070]=30'd260631016;
array2[7071]=30'd228181405;
array2[7072]=30'd265928088;
array2[7073]=30'd281654691;
array2[7074]=30'd269069720;
array2[7075]=30'd221916546;
array2[7076]=30'd230307208;
array2[7077]=30'd227165569;
array2[7078]=30'd231362949;
array2[7079]=30'd231362949;
array2[7080]=30'd231362949;
array2[7081]=30'd231362949;
array2[7082]=30'd231362949;
array2[7083]=30'd234504581;
array2[7084]=30'd234504581;
array2[7085]=30'd231364996;
array2[7086]=30'd230317442;
array2[7087]=30'd231364996;
array2[7088]=30'd229266819;
array2[7089]=30'd231362949;
array2[7090]=30'd229266819;
array2[7091]=30'd231362949;
array2[7092]=30'd229266819;
array2[7093]=30'd234504581;
array2[7094]=30'd231362949;
array2[7095]=30'd231362949;
array2[7096]=30'd227165569;
array2[7097]=30'd231362949;
array2[7098]=30'd228216193;
array2[7099]=30'd231362949;
array2[7100]=30'd234504581;
array2[7101]=30'd231362949;
array2[7102]=30'd228216193;
array2[7103]=30'd231362949;
array2[7104]=30'd193577377;
array2[7105]=30'd234504581;
array2[7106]=30'd227165569;
array2[7107]=30'd228216193;
array2[7108]=30'd230317442;
array2[7109]=30'd231362949;
array2[7110]=30'd229266819;
array2[7111]=30'd230317442;
array2[7112]=30'd232417668;
array2[7113]=30'd229266819;
array2[7114]=30'd231362949;
array2[7115]=30'd232417668;
array2[7116]=30'd229266819;
array2[7117]=30'd231362949;
array2[7118]=30'd229266819;
array2[7119]=30'd231359873;
array2[7120]=30'd229266819;
array2[7121]=30'd230317442;
array2[7122]=30'd231362949;
array2[7123]=30'd229266819;
array2[7124]=30'd231364996;
array2[7125]=30'd231362949;
array2[7126]=30'd231362949;
array2[7127]=30'd236604812;
array2[7128]=30'd231362949;
array2[7129]=30'd231362949;
array2[7130]=30'd234504581;
array2[7131]=30'd234504581;
array2[7132]=30'd304706973;
array2[7133]=30'd295249323;
array2[7134]=30'd271165847;
array2[7135]=30'd262793620;
array2[7136]=30'd248105365;
array2[7137]=30'd240774546;
array2[7138]=30'd212454818;
array2[7139]=30'd218607140;
array2[7140]=30'd331763301;
array2[7141]=30'd265736724;
array2[7142]=30'd193577377;
array2[7143]=30'd213516691;
array2[7144]=30'd213516691;
array2[7145]=30'd228216193;
array2[7146]=30'd231364996;
array2[7147]=30'd231362949;
array2[7148]=30'd229266819;
array2[7149]=30'd231364996;
array2[7150]=30'd236604812;
array2[7151]=30'd256519562;
array2[7152]=30'd220861839;
array2[7153]=30'd212454818;
array2[7154]=30'd212454818;
array2[7155]=30'd190356956;
array2[7156]=30'd124307934;
array2[7157]=30'd106464746;
array2[7158]=30'd124307934;
array2[7159]=30'd131612152;
array2[7160]=30'd407216718;
array2[7161]=30'd299264555;
array2[7162]=30'd407216718;
array2[7163]=30'd604201637;
array2[7164]=30'd601041592;
array2[7165]=30'd560184961;
array2[7166]=30'd407216718;
array2[7167]=30'd319215128;
array2[7168]=30'd254365107;
array2[7169]=30'd271165847;
array2[7170]=30'd257539480;
array2[7171]=30'd265928088;
array2[7172]=30'd265928088;
array2[7173]=30'd227159434;
array2[7174]=30'd262793620;
array2[7175]=30'd262793620;
array2[7176]=30'd262793620;
array2[7177]=30'd234499470;
array2[7178]=30'd231362949;
array2[7179]=30'd231362949;
array2[7180]=30'd228216193;
array2[7181]=30'd230317442;
array2[7182]=30'd229266819;
array2[7183]=30'd231362949;
array2[7184]=30'd229266819;
array2[7185]=30'd229266819;
array2[7186]=30'd229266819;
array2[7187]=30'd231362949;
array2[7188]=30'd229266819;
array2[7189]=30'd231362949;
array2[7190]=30'd229266819;
array2[7191]=30'd229266819;
array2[7192]=30'd231362949;
array2[7193]=30'd231362949;
array2[7194]=30'd229266819;
array2[7195]=30'd230317442;
array2[7196]=30'd231362949;
array2[7197]=30'd228216193;
array2[7198]=30'd231362949;
array2[7199]=30'd230317442;
array2[7200]=30'd193577377;
array2[7201]=30'd234504581;
array2[7202]=30'd227165569;
array2[7203]=30'd228216193;
array2[7204]=30'd229266819;
array2[7205]=30'd229266819;
array2[7206]=30'd229266819;
array2[7207]=30'd229266819;
array2[7208]=30'd230317442;
array2[7209]=30'd229266819;
array2[7210]=30'd231362949;
array2[7211]=30'd229270912;
array2[7212]=30'd228216193;
array2[7213]=30'd231362949;
array2[7214]=30'd229266819;
array2[7215]=30'd231359873;
array2[7216]=30'd229266819;
array2[7217]=30'd229266819;
array2[7218]=30'd231362949;
array2[7219]=30'd229266819;
array2[7220]=30'd229266819;
array2[7221]=30'd234504581;
array2[7222]=30'd234504581;
array2[7223]=30'd231362949;
array2[7224]=30'd231362949;
array2[7225]=30'd227165569;
array2[7226]=30'd231362949;
array2[7227]=30'd227165569;
array2[7228]=30'd271165847;
array2[7229]=30'd304706973;
array2[7230]=30'd295249323;
array2[7231]=30'd312021416;
array2[7232]=30'd304706973;
array2[7233]=30'd271165847;
array2[7234]=30'd212454818;
array2[7235]=30'd159912438;
array2[7236]=30'd299264555;
array2[7237]=30'd331763301;
array2[7238]=30'd299264555;
array2[7239]=30'd299264555;
array2[7240]=30'd218607140;
array2[7241]=30'd228181405;
array2[7242]=30'd228216193;
array2[7243]=30'd228212100;
array2[7244]=30'd231359873;
array2[7245]=30'd229266819;
array2[7246]=30'd230307208;
array2[7247]=30'd207191473;
array2[7248]=30'd260631016;
array2[7249]=30'd265736724;
array2[7250]=30'd299264555;
array2[7251]=30'd295074390;
array2[7252]=30'd347490866;
array2[7253]=30'd124307934;
array2[7254]=30'd106464746;
array2[7255]=30'd124307934;
array2[7256]=30'd645112409;
array2[7257]=30'd646130287;
array2[7258]=30'd631447172;
array2[7259]=30'd606320275;
array2[7260]=30'd606320275;
array2[7261]=30'd604201637;
array2[7262]=30'd604201637;
array2[7263]=30'd560184961;
array2[7264]=30'd383147560;
array2[7265]=30'd260631016;
array2[7266]=30'd254365107;
array2[7267]=30'd280599950;
array2[7268]=30'd304706973;
array2[7269]=30'd295249323;
array2[7270]=30'd304706973;
array2[7271]=30'd304706973;
array2[7272]=30'd312021416;
array2[7273]=30'd271165847;
array2[7274]=30'd257539480;
array2[7275]=30'd221916546;
array2[7276]=30'd230307208;
array2[7277]=30'd231362949;
array2[7278]=30'd231362949;
array2[7279]=30'd231362949;
array2[7280]=30'd231362949;
array2[7281]=30'd231362949;
array2[7282]=30'd231362949;
array2[7283]=30'd231362949;
array2[7284]=30'd229266819;
array2[7285]=30'd231362949;
array2[7286]=30'd229266819;
array2[7287]=30'd229266819;
array2[7288]=30'd231362949;
array2[7289]=30'd231362949;
array2[7290]=30'd229266819;
array2[7291]=30'd231362949;
array2[7292]=30'd231362949;
array2[7293]=30'd231364996;
array2[7294]=30'd231364996;
array2[7295]=30'd229266819;
array2[7296]=30'd193577377;
array2[7297]=30'd234504581;
array2[7298]=30'd227165569;
array2[7299]=30'd234504581;
array2[7300]=30'd232392085;
array2[7301]=30'd232392085;
array2[7302]=30'd232392085;
array2[7303]=30'd232392085;
array2[7304]=30'd227159434;
array2[7305]=30'd232392085;
array2[7306]=30'd232392085;
array2[7307]=30'd227159434;
array2[7308]=30'd232392085;
array2[7309]=30'd232392085;
array2[7310]=30'd232392085;
array2[7311]=30'd232392085;
array2[7312]=30'd225072515;
array2[7313]=30'd231364996;
array2[7314]=30'd231362949;
array2[7315]=30'd231362949;
array2[7316]=30'd229270912;
array2[7317]=30'd228216193;
array2[7318]=30'd231364996;
array2[7319]=30'd231364996;
array2[7320]=30'd234504581;
array2[7321]=30'd229266819;
array2[7322]=30'd231364996;
array2[7323]=30'd234499470;
array2[7324]=30'd257539480;
array2[7325]=30'd248105365;
array2[7326]=30'd228181405;
array2[7327]=30'd248105365;
array2[7328]=30'd267996623;
array2[7329]=30'd295249323;
array2[7330]=30'd267996623;
array2[7331]=30'd207191473;
array2[7332]=30'd190356956;
array2[7333]=30'd249001484;
array2[7334]=30'd265736724;
array2[7335]=30'd265736724;
array2[7336]=30'd299264555;
array2[7337]=30'd195647926;
array2[7338]=30'd227165569;
array2[7339]=30'd230307208;
array2[7340]=30'd231362949;
array2[7341]=30'd227159434;
array2[7342]=30'd260631016;
array2[7343]=30'd506770009;
array2[7344]=30'd449120871;
array2[7345]=30'd357913199;
array2[7346]=30'd357913199;
array2[7347]=30'd434416250;
array2[7348]=30'd606320275;
array2[7349]=30'd449120871;
array2[7350]=30'd299264555;
array2[7351]=30'd124307934;
array2[7352]=30'd646130287;
array2[7353]=30'd764529268;
array2[7354]=30'd768729747;
array2[7355]=30'd768729747;
array2[7356]=30'd672348794;
array2[7357]=30'd560184961;
array2[7358]=30'd560184961;
array2[7359]=30'd604201637;
array2[7360]=30'd539218630;
array2[7361]=30'd481587821;
array2[7362]=30'd319215128;
array2[7363]=30'd254365107;
array2[7364]=30'd304706973;
array2[7365]=30'd312021416;
array2[7366]=30'd295249323;
array2[7367]=30'd304706973;
array2[7368]=30'd312021416;
array2[7369]=30'd304706973;
array2[7370]=30'd280599950;
array2[7371]=30'd248105365;
array2[7372]=30'd238691720;
array2[7373]=30'd227165569;
array2[7374]=30'd231359873;
array2[7375]=30'd231362949;
array2[7376]=30'd231364996;
array2[7377]=30'd231362949;
array2[7378]=30'd231362949;
array2[7379]=30'd231362949;
array2[7380]=30'd231362949;
array2[7381]=30'd231362949;
array2[7382]=30'd228216193;
array2[7383]=30'd229266819;
array2[7384]=30'd228216193;
array2[7385]=30'd231362949;
array2[7386]=30'd229266819;
array2[7387]=30'd231362949;
array2[7388]=30'd234504581;
array2[7389]=30'd227165569;
array2[7390]=30'd229266819;
array2[7391]=30'd234504581;
array2[7392]=30'd260631016;
array2[7393]=30'd267996623;
array2[7394]=30'd280568333;
array2[7395]=30'd284737060;
array2[7396]=30'd390446940;
array2[7397]=30'd461700935;
array2[7398]=30'd461700935;
array2[7399]=30'd461700935;
array2[7400]=30'd461700935;
array2[7401]=30'd461700935;
array2[7402]=30'd461700935;
array2[7403]=30'd461700935;
array2[7404]=30'd461700935;
array2[7405]=30'd461700935;
array2[7406]=30'd461700935;
array2[7407]=30'd328674981;
array2[7408]=30'd280568333;
array2[7409]=30'd280568333;
array2[7410]=30'd280568333;
array2[7411]=30'd280568333;
array2[7412]=30'd280568333;
array2[7413]=30'd280568333;
array2[7414]=30'd280568333;
array2[7415]=30'd280568333;
array2[7416]=30'd280568333;
array2[7417]=30'd280568333;
array2[7418]=30'd280568333;
array2[7419]=30'd357996288;
array2[7420]=30'd461700935;
array2[7421]=30'd461700935;
array2[7422]=30'd461700935;
array2[7423]=30'd461700935;
array2[7424]=30'd461700935;
array2[7425]=30'd461700935;
array2[7426]=30'd461700935;
array2[7427]=30'd461700935;
array2[7428]=30'd390446940;
array2[7429]=30'd451191548;
array2[7430]=30'd357996288;
array2[7431]=30'd178773498;
array2[7432]=30'd295074390;
array2[7433]=30'd218607140;
array2[7434]=30'd195647926;
array2[7435]=30'd267996623;
array2[7436]=30'd280568333;
array2[7437]=30'd260631016;
array2[7438]=30'd560184961;
array2[7439]=30'd713179821;
array2[7440]=30'd565444213;
array2[7441]=30'd357913199;
array2[7442]=30'd357913199;
array2[7443]=30'd449120871;
array2[7444]=30'd711090860;
array2[7445]=30'd678602388;
array2[7446]=30'd434416250;
array2[7447]=30'd218607140;
array2[7448]=30'd407216718;
array2[7449]=30'd711090860;
array2[7450]=30'd819020415;
array2[7451]=30'd828452495;
array2[7452]=30'd819020415;
array2[7453]=30'd727851632;
array2[7454]=30'd677571193;
array2[7455]=30'd560184961;
array2[7456]=30'd560184961;
array2[7457]=30'd518272648;
array2[7458]=30'd483727963;
array2[7459]=30'd319215128;
array2[7460]=30'd260631016;
array2[7461]=30'd260631016;
array2[7462]=30'd312021416;
array2[7463]=30'd312021416;
array2[7464]=30'd312021416;
array2[7465]=30'd304706973;
array2[7466]=30'd304706973;
array2[7467]=30'd312021416;
array2[7468]=30'd269069720;
array2[7469]=30'd230307208;
array2[7470]=30'd231359873;
array2[7471]=30'd231362949;
array2[7472]=30'd231364996;
array2[7473]=30'd231362949;
array2[7474]=30'd231362949;
array2[7475]=30'd231362949;
array2[7476]=30'd229266819;
array2[7477]=30'd231362949;
array2[7478]=30'd231359873;
array2[7479]=30'd229266819;
array2[7480]=30'd228216193;
array2[7481]=30'd229266819;
array2[7482]=30'd229266819;
array2[7483]=30'd231362949;
array2[7484]=30'd234504581;
array2[7485]=30'd227165569;
array2[7486]=30'd229266819;
array2[7487]=30'd231362949;
array2[7488]=30'd390446940;
array2[7489]=30'd409311115;
array2[7490]=30'd409311115;
array2[7491]=30'd409311115;
array2[7492]=30'd429185963;
array2[7493]=30'd426044336;
array2[7494]=30'd426044336;
array2[7495]=30'd423950257;
array2[7496]=30'd423950257;
array2[7497]=30'd423950257;
array2[7498]=30'd423950257;
array2[7499]=30'd426044336;
array2[7500]=30'd423950257;
array2[7501]=30'd423950257;
array2[7502]=30'd429185963;
array2[7503]=30'd429185963;
array2[7504]=30'd409311115;
array2[7505]=30'd409311115;
array2[7506]=30'd409311115;
array2[7507]=30'd409311115;
array2[7508]=30'd409311115;
array2[7509]=30'd409311115;
array2[7510]=30'd409311115;
array2[7511]=30'd409311115;
array2[7512]=30'd409311115;
array2[7513]=30'd409311115;
array2[7514]=30'd409311115;
array2[7515]=30'd429185963;
array2[7516]=30'd426044336;
array2[7517]=30'd423950257;
array2[7518]=30'd423950257;
array2[7519]=30'd423950257;
array2[7520]=30'd423950257;
array2[7521]=30'd426044336;
array2[7522]=30'd426044336;
array2[7523]=30'd426044336;
array2[7524]=30'd423950257;
array2[7525]=30'd423950257;
array2[7526]=30'd409311115;
array2[7527]=30'd287786593;
array2[7528]=30'd295074390;
array2[7529]=30'd357913199;
array2[7530]=30'd339090072;
array2[7531]=30'd218607140;
array2[7532]=30'd299264555;
array2[7533]=30'd604201637;
array2[7534]=30'd770812573;
array2[7535]=30'd819020415;
array2[7536]=30'd645112409;
array2[7537]=30'd357913199;
array2[7538]=30'd434416250;
array2[7539]=30'd481587821;
array2[7540]=30'd768729747;
array2[7541]=30'd768729747;
array2[7542]=30'd565444213;
array2[7543]=30'd375721588;
array2[7544]=30'd265736724;
array2[7545]=30'd566515308;
array2[7546]=30'd713179821;
array2[7547]=30'd819020415;
array2[7548]=30'd851505800;
array2[7549]=30'd828452495;
array2[7550]=30'd828452495;
array2[7551]=30'd768729747;
array2[7552]=30'd678602388;
array2[7553]=30'd604201637;
array2[7554]=30'd768729747;
array2[7555]=30'd790726247;
array2[7556]=30'd764529268;
array2[7557]=30'd678602388;
array2[7558]=30'd281508345;
array2[7559]=30'd249001484;
array2[7560]=30'd254365107;
array2[7561]=30'd304706973;
array2[7562]=30'd295249323;
array2[7563]=30'd304706973;
array2[7564]=30'd280599950;
array2[7565]=30'd227159434;
array2[7566]=30'd227165569;
array2[7567]=30'd231362949;
array2[7568]=30'd231362949;
array2[7569]=30'd231362949;
array2[7570]=30'd230317442;
array2[7571]=30'd230317442;
array2[7572]=30'd229266819;
array2[7573]=30'd231362949;
array2[7574]=30'd229266819;
array2[7575]=30'd229266819;
array2[7576]=30'd229266819;
array2[7577]=30'd230317442;
array2[7578]=30'd229266819;
array2[7579]=30'd231362949;
array2[7580]=30'd231362949;
array2[7581]=30'd229266819;
array2[7582]=30'd231362949;
array2[7583]=30'd231364996;
array2[7584]=30'd390446940;
array2[7585]=30'd426044336;
array2[7586]=30'd426044336;
array2[7587]=30'd423950257;
array2[7588]=30'd423950257;
array2[7589]=30'd426044336;
array2[7590]=30'd426044336;
array2[7591]=30'd423950257;
array2[7592]=30'd423950257;
array2[7593]=30'd423950257;
array2[7594]=30'd426044336;
array2[7595]=30'd426044336;
array2[7596]=30'd423950257;
array2[7597]=30'd426044336;
array2[7598]=30'd426044336;
array2[7599]=30'd426044336;
array2[7600]=30'd426044336;
array2[7601]=30'd423950257;
array2[7602]=30'd423950257;
array2[7603]=30'd423950257;
array2[7604]=30'd423950257;
array2[7605]=30'd423950257;
array2[7606]=30'd426044336;
array2[7607]=30'd426044336;
array2[7608]=30'd426044336;
array2[7609]=30'd423950257;
array2[7610]=30'd423950257;
array2[7611]=30'd426044336;
array2[7612]=30'd426044336;
array2[7613]=30'd426044336;
array2[7614]=30'd426044336;
array2[7615]=30'd423950257;
array2[7616]=30'd426044336;
array2[7617]=30'd426044336;
array2[7618]=30'd426044336;
array2[7619]=30'd426044336;
array2[7620]=30'd426044336;
array2[7621]=30'd426044336;
array2[7622]=30'd426044336;
array2[7623]=30'd429185963;
array2[7624]=30'd390446940;
array2[7625]=30'd287786593;
array2[7626]=30'd218607140;
array2[7627]=30'd295074390;
array2[7628]=30'd601041592;
array2[7629]=30'd770816666;
array2[7630]=30'd790726247;
array2[7631]=30'd805398138;
array2[7632]=30'd768729747;
array2[7633]=30'd560184961;
array2[7634]=30'd449120871;
array2[7635]=30'd518272648;
array2[7636]=30'd805398138;
array2[7637]=30'd819020415;
array2[7638]=30'd565444213;
array2[7639]=30'd450208341;
array2[7640]=30'd380968597;
array2[7641]=30'd606320275;
array2[7642]=30'd566515308;
array2[7643]=30'd606320275;
array2[7644]=30'd768729747;
array2[7645]=30'd819020415;
array2[7646]=30'd828452495;
array2[7647]=30'd851505800;
array2[7648]=30'd851505800;
array2[7649]=30'd828452495;
array2[7650]=30'd851505800;
array2[7651]=30'd858839683;
array2[7652]=30'd858839683;
array2[7653]=30'd851505800;
array2[7654]=30'd819020415;
array2[7655]=30'd768729747;
array2[7656]=30'd506770009;
array2[7657]=30'd265736724;
array2[7658]=30'd260631016;
array2[7659]=30'd271165847;
array2[7660]=30'd280599950;
array2[7661]=30'd265928088;
array2[7662]=30'd238691720;
array2[7663]=30'd231362949;
array2[7664]=30'd230317442;
array2[7665]=30'd231364996;
array2[7666]=30'd231364996;
array2[7667]=30'd231362949;
array2[7668]=30'd229266819;
array2[7669]=30'd231362949;
array2[7670]=30'd229266819;
array2[7671]=30'd229266819;
array2[7672]=30'd229266819;
array2[7673]=30'd228216193;
array2[7674]=30'd229266819;
array2[7675]=30'd231362949;
array2[7676]=30'd231359873;
array2[7677]=30'd231362949;
array2[7678]=30'd227165569;
array2[7679]=30'd231362949;
array2[7680]=30'd390446940;
array2[7681]=30'd426044336;
array2[7682]=30'd435467177;
array2[7683]=30'd435467177;
array2[7684]=30'd635645720;
array2[7685]=30'd672324351;
array2[7686]=30'd672324351;
array2[7687]=30'd672324351;
array2[7688]=30'd672324351;
array2[7689]=30'd672324351;
array2[7690]=30'd672324351;
array2[7691]=30'd672324351;
array2[7692]=30'd672324351;
array2[7693]=30'd672324351;
array2[7694]=30'd672324351;
array2[7695]=30'd493111164;
array2[7696]=30'd426044336;
array2[7697]=30'd426044336;
array2[7698]=30'd426044336;
array2[7699]=30'd426044336;
array2[7700]=30'd426044336;
array2[7701]=30'd426044336;
array2[7702]=30'd426044336;
array2[7703]=30'd426044336;
array2[7704]=30'd426044336;
array2[7705]=30'd426044336;
array2[7706]=30'd435467177;
array2[7707]=30'd582196031;
array2[7708]=30'd672324351;
array2[7709]=30'd672324351;
array2[7710]=30'd672324351;
array2[7711]=30'd672324351;
array2[7712]=30'd672324351;
array2[7713]=30'd672324351;
array2[7714]=30'd672324351;
array2[7715]=30'd672324351;
array2[7716]=30'd672324351;
array2[7717]=30'd672324351;
array2[7718]=30'd582196031;
array2[7719]=30'd426044336;
array2[7720]=30'd429185963;
array2[7721]=30'd429185963;
array2[7722]=30'd395649781;
array2[7723]=30'd339090072;
array2[7724]=30'd711090860;
array2[7725]=30'd805398138;
array2[7726]=30'd805398138;
array2[7727]=30'd805398138;
array2[7728]=30'd828452495;
array2[7729]=30'd678602388;
array2[7730]=30'd434416250;
array2[7731]=30'd506770009;
array2[7732]=30'd823228019;
array2[7733]=30'd819020415;
array2[7734]=30'd560184961;
array2[7735]=30'd434416250;
array2[7736]=30'd560184961;
array2[7737]=30'd768729747;
array2[7738]=30'd770812573;
array2[7739]=30'd678602388;
array2[7740]=30'd560184961;
array2[7741]=30'd672348794;
array2[7742]=30'd727851632;
array2[7743]=30'd819020415;
array2[7744]=30'd851505800;
array2[7745]=30'd851505800;
array2[7746]=30'd858839683;
array2[7747]=30'd858839683;
array2[7748]=30'd858839683;
array2[7749]=30'd865130113;
array2[7750]=30'd858839683;
array2[7751]=30'd851505800;
array2[7752]=30'd851505800;
array2[7753]=30'd768729747;
array2[7754]=30'd450208341;
array2[7755]=30'd254365107;
array2[7756]=30'd280599950;
array2[7757]=30'd271165847;
array2[7758]=30'd227165569;
array2[7759]=30'd231359873;
array2[7760]=30'd231364996;
array2[7761]=30'd230317442;
array2[7762]=30'd231362949;
array2[7763]=30'd231359873;
array2[7764]=30'd231362949;
array2[7765]=30'd231362949;
array2[7766]=30'd231362949;
array2[7767]=30'd231362949;
array2[7768]=30'd228216193;
array2[7769]=30'd231362949;
array2[7770]=30'd231362949;
array2[7771]=30'd231362949;
array2[7772]=30'd231362949;
array2[7773]=30'd228216193;
array2[7774]=30'd234504581;
array2[7775]=30'd231359873;
array2[7776]=30'd601041592;
array2[7777]=30'd672324351;
array2[7778]=30'd672324351;
array2[7779]=30'd718417640;
array2[7780]=30'd718417640;
array2[7781]=30'd728897252;
array2[7782]=30'd728897252;
array2[7783]=30'd728897252;
array2[7784]=30'd728897252;
array2[7785]=30'd728897252;
array2[7786]=30'd728897252;
array2[7787]=30'd728897252;
array2[7788]=30'd728897252;
array2[7789]=30'd728897252;
array2[7790]=30'd728897252;
array2[7791]=30'd718417640;
array2[7792]=30'd672324351;
array2[7793]=30'd672324351;
array2[7794]=30'd672324351;
array2[7795]=30'd672324351;
array2[7796]=30'd672324351;
array2[7797]=30'd672324351;
array2[7798]=30'd672324351;
array2[7799]=30'd672324351;
array2[7800]=30'd672324351;
array2[7801]=30'd718417640;
array2[7802]=30'd672324351;
array2[7803]=30'd718417640;
array2[7804]=30'd718417640;
array2[7805]=30'd728897252;
array2[7806]=30'd728897252;
array2[7807]=30'd718417640;
array2[7808]=30'd718417640;
array2[7809]=30'd718417640;
array2[7810]=30'd718417640;
array2[7811]=30'd718417640;
array2[7812]=30'd718417640;
array2[7813]=30'd718417640;
array2[7814]=30'd718417640;
array2[7815]=30'd718417640;
array2[7816]=30'd718417640;
array2[7817]=30'd672324351;
array2[7818]=30'd539218630;
array2[7819]=30'd606320275;
array2[7820]=30'd770816666;
array2[7821]=30'd805398138;
array2[7822]=30'd823228019;
array2[7823]=30'd805398138;
array2[7824]=30'd828452495;
array2[7825]=30'd799112870;
array2[7826]=30'd672348794;
array2[7827]=30'd678604396;
array2[7828]=30'd851505800;
array2[7829]=30'd828452495;
array2[7830]=30'd645112409;
array2[7831]=30'd434416250;
array2[7832]=30'd711090860;
array2[7833]=30'd828452495;
array2[7834]=30'd851505800;
array2[7835]=30'd828452495;
array2[7836]=30'd768729747;
array2[7837]=30'd631447172;
array2[7838]=30'd565444213;
array2[7839]=30'd678602388;
array2[7840]=30'd768729747;
array2[7841]=30'd851505800;
array2[7842]=30'd851505800;
array2[7843]=30'd858839683;
array2[7844]=30'd858839683;
array2[7845]=30'd858839683;
array2[7846]=30'd858839683;
array2[7847]=30'd858839683;
array2[7848]=30'd858839683;
array2[7849]=30'd851505800;
array2[7850]=30'd727851632;
array2[7851]=30'd190356956;
array2[7852]=30'd280599950;
array2[7853]=30'd280599950;
array2[7854]=30'd227165569;
array2[7855]=30'd231362949;
array2[7856]=30'd231362949;
array2[7857]=30'd231359873;
array2[7858]=30'd231362949;
array2[7859]=30'd231359873;
array2[7860]=30'd231359873;
array2[7861]=30'd231362949;
array2[7862]=30'd228216193;
array2[7863]=30'd231362949;
array2[7864]=30'd231362949;
array2[7865]=30'd231362949;
array2[7866]=30'd231362949;
array2[7867]=30'd230317442;
array2[7868]=30'd231362949;
array2[7869]=30'd230317442;
array2[7870]=30'd231362949;
array2[7871]=30'd231362949;
array2[7872]=30'd646169309;
array2[7873]=30'd718417640;
array2[7874]=30'd728897252;
array2[7875]=30'd728897252;
array2[7876]=30'd728897252;
array2[7877]=30'd728897252;
array2[7878]=30'd728897252;
array2[7879]=30'd728897252;
array2[7880]=30'd728897252;
array2[7881]=30'd728897252;
array2[7882]=30'd728897252;
array2[7883]=30'd728897252;
array2[7884]=30'd728897252;
array2[7885]=30'd728897252;
array2[7886]=30'd728897252;
array2[7887]=30'd728897252;
array2[7888]=30'd728897252;
array2[7889]=30'd728897252;
array2[7890]=30'd728897252;
array2[7891]=30'd728897252;
array2[7892]=30'd728897252;
array2[7893]=30'd728897252;
array2[7894]=30'd728897252;
array2[7895]=30'd728897252;
array2[7896]=30'd728897252;
array2[7897]=30'd728897252;
array2[7898]=30'd728897252;
array2[7899]=30'd728897252;
array2[7900]=30'd728897252;
array2[7901]=30'd728897252;
array2[7902]=30'd728897252;
array2[7903]=30'd728897252;
array2[7904]=30'd728897252;
array2[7905]=30'd728897252;
array2[7906]=30'd728897252;
array2[7907]=30'd718417640;
array2[7908]=30'd718417640;
array2[7909]=30'd718417640;
array2[7910]=30'd718417640;
array2[7911]=30'd728897252;
array2[7912]=30'd728897252;
array2[7913]=30'd601041592;
array2[7914]=30'd481587821;
array2[7915]=30'd764529268;
array2[7916]=30'd828452495;
array2[7917]=30'd828452495;
array2[7918]=30'd823228019;
array2[7919]=30'd823228019;
array2[7920]=30'd828452495;
array2[7921]=30'd851505800;
array2[7922]=30'd851505800;
array2[7923]=30'd858839683;
array2[7924]=30'd858839683;
array2[7925]=30'd851505800;
array2[7926]=30'd764529268;
array2[7927]=30'd727851632;
array2[7928]=30'd819020415;
array2[7929]=30'd851505800;
array2[7930]=30'd858839683;
array2[7931]=30'd858839683;
array2[7932]=30'd858839683;
array2[7933]=30'd828452495;
array2[7934]=30'd799112870;
array2[7935]=30'd764529268;
array2[7936]=30'd805398138;
array2[7937]=30'd851505800;
array2[7938]=30'd858839683;
array2[7939]=30'd858839683;
array2[7940]=30'd858839683;
array2[7941]=30'd858839683;
array2[7942]=30'd858839683;
array2[7943]=30'd851505800;
array2[7944]=30'd858839683;
array2[7945]=30'd858839683;
array2[7946]=30'd770816666;
array2[7947]=30'd506770009;
array2[7948]=30'd260631016;
array2[7949]=30'd271165847;
array2[7950]=30'd232392085;
array2[7951]=30'd232417668;
array2[7952]=30'd231364996;
array2[7953]=30'd229266819;
array2[7954]=30'd229266819;
array2[7955]=30'd229266819;
array2[7956]=30'd231362949;
array2[7957]=30'd231362949;
array2[7958]=30'd231362949;
array2[7959]=30'd230317442;
array2[7960]=30'd231362949;
array2[7961]=30'd230317442;
array2[7962]=30'd231362949;
array2[7963]=30'd231362949;
array2[7964]=30'd229266819;
array2[7965]=30'd231364996;
array2[7966]=30'd229266819;
array2[7967]=30'd229266819;
array2[7968]=30'd678602388;
array2[7969]=30'd728897252;
array2[7970]=30'd728897252;
array2[7971]=30'd758240964;
array2[7972]=30'd828452495;
array2[7973]=30'd858839683;
array2[7974]=30'd865130113;
array2[7975]=30'd858839683;
array2[7976]=30'd865130113;
array2[7977]=30'd858839683;
array2[7978]=30'd865130113;
array2[7979]=30'd865130113;
array2[7980]=30'd858839683;
array2[7981]=30'd865130113;
array2[7982]=30'd865130113;
array2[7983]=30'd799112870;
array2[7984]=30'd728897252;
array2[7985]=30'd728897252;
array2[7986]=30'd728897252;
array2[7987]=30'd728897252;
array2[7988]=30'd728897252;
array2[7989]=30'd728897252;
array2[7990]=30'd728897252;
array2[7991]=30'd728897252;
array2[7992]=30'd728897252;
array2[7993]=30'd728897252;
array2[7994]=30'd728897252;
array2[7995]=30'd828452495;
array2[7996]=30'd858839683;
array2[7997]=30'd865130113;
array2[7998]=30'd865130113;
array2[7999]=30'd865130113;
array2[8000]=30'd858839683;
array2[8001]=30'd865130113;
array2[8002]=30'd865130113;
array2[8003]=30'd851505800;
array2[8004]=30'd770812573;
array2[8005]=30'd805398138;
array2[8006]=30'd770816666;
array2[8007]=30'd732038833;
array2[8008]=30'd718417640;
array2[8009]=30'd606320275;
array2[8010]=30'd506770009;
array2[8011]=30'd851505800;
array2[8012]=30'd828452495;
array2[8013]=30'd858839683;
array2[8014]=30'd828452495;
array2[8015]=30'd805398138;
array2[8016]=30'd819020415;
array2[8017]=30'd828452495;
array2[8018]=30'd851505800;
array2[8019]=30'd851505800;
array2[8020]=30'd858839683;
array2[8021]=30'd858839683;
array2[8022]=30'd819020415;
array2[8023]=30'd828452495;
array2[8024]=30'd858839683;
array2[8025]=30'd851505800;
array2[8026]=30'd858839683;
array2[8027]=30'd858839683;
array2[8028]=30'd858839683;
array2[8029]=30'd858839683;
array2[8030]=30'd858839683;
array2[8031]=30'd851505800;
array2[8032]=30'd858839683;
array2[8033]=30'd858839683;
array2[8034]=30'd858839683;
array2[8035]=30'd858839683;
array2[8036]=30'd858839683;
array2[8037]=30'd851505800;
array2[8038]=30'd828452495;
array2[8039]=30'd851505800;
array2[8040]=30'd851505800;
array2[8041]=30'd858839683;
array2[8042]=30'd828452495;
array2[8043]=30'd678602388;
array2[8044]=30'd281508345;
array2[8045]=30'd280599950;
array2[8046]=30'd240774546;
array2[8047]=30'd227165569;
array2[8048]=30'd229266819;
array2[8049]=30'd231362949;
array2[8050]=30'd234504581;
array2[8051]=30'd228216193;
array2[8052]=30'd231364996;
array2[8053]=30'd231362949;
array2[8054]=30'd231362949;
array2[8055]=30'd231362949;
array2[8056]=30'd231362949;
array2[8057]=30'd231362949;
array2[8058]=30'd231362949;
array2[8059]=30'd231362949;
array2[8060]=30'd228216193;
array2[8061]=30'd229266819;
array2[8062]=30'd231362949;
array2[8063]=30'd231362949;
array2[8064]=30'd764529268;
array2[8065]=30'd865130113;
array2[8066]=30'd858839683;
array2[8067]=30'd865130113;
array2[8068]=30'd906004072;
array2[8069]=30'd906004072;
array2[8070]=30'd906004072;
array2[8071]=30'd906004072;
array2[8072]=30'd906004072;
array2[8073]=30'd906004072;
array2[8074]=30'd906004072;
array2[8075]=30'd906004072;
array2[8076]=30'd906004072;
array2[8077]=30'd906004072;
array2[8078]=30'd906004072;
array2[8079]=30'd906004072;
array2[8080]=30'd865130113;
array2[8081]=30'd865130113;
array2[8082]=30'd865130113;
array2[8083]=30'd865130113;
array2[8084]=30'd865130113;
array2[8085]=30'd865130113;
array2[8086]=30'd865130113;
array2[8087]=30'd865130113;
array2[8088]=30'd865130113;
array2[8089]=30'd865130113;
array2[8090]=30'd851505800;
array2[8091]=30'd906004072;
array2[8092]=30'd906004072;
array2[8093]=30'd906004072;
array2[8094]=30'd906004072;
array2[8095]=30'd906004072;
array2[8096]=30'd906004072;
array2[8097]=30'd906004072;
array2[8098]=30'd906004072;
array2[8099]=30'd906004072;
array2[8100]=30'd823228019;
array2[8101]=30'd858839683;
array2[8102]=30'd823228019;
array2[8103]=30'd805398138;
array2[8104]=30'd819020415;
array2[8105]=30'd678604396;
array2[8106]=30'd538207812;
array2[8107]=30'd858839683;
array2[8108]=30'd851505800;
array2[8109]=30'd858839683;
array2[8110]=30'd858839683;
array2[8111]=30'd819020415;
array2[8112]=30'd819020415;
array2[8113]=30'd828452495;
array2[8114]=30'd858839683;
array2[8115]=30'd858839683;
array2[8116]=30'd858839683;
array2[8117]=30'd858839683;
array2[8118]=30'd858839683;
array2[8119]=30'd858839683;
array2[8120]=30'd858839683;
array2[8121]=30'd858839683;
array2[8122]=30'd851505800;
array2[8123]=30'd858839683;
array2[8124]=30'd851505800;
array2[8125]=30'd858839683;
array2[8126]=30'd858839683;
array2[8127]=30'd858839683;
array2[8128]=30'd858839683;
array2[8129]=30'd858839683;
array2[8130]=30'd865130113;
array2[8131]=30'd851505800;
array2[8132]=30'd858839683;
array2[8133]=30'd828452495;
array2[8134]=30'd828452495;
array2[8135]=30'd819020415;
array2[8136]=30'd805398138;
array2[8137]=30'd805398138;
array2[8138]=30'd851505800;
array2[8139]=30'd762499681;
array2[8140]=30'd281508345;
array2[8141]=30'd304706973;
array2[8142]=30'd295249323;
array2[8143]=30'd240774546;
array2[8144]=30'd238691720;
array2[8145]=30'd230307208;
array2[8146]=30'd225072515;
array2[8147]=30'd229266819;
array2[8148]=30'd231364996;
array2[8149]=30'd228216193;
array2[8150]=30'd231362949;
array2[8151]=30'd230317442;
array2[8152]=30'd231364996;
array2[8153]=30'd231362949;
array2[8154]=30'd231362949;
array2[8155]=30'd231362949;
array2[8156]=30'd231362949;
array2[8157]=30'd227165569;
array2[8158]=30'd228216193;
array2[8159]=30'd227165569;
array2[8160]=30'd790726247;
array2[8161]=30'd906004072;
array2[8162]=30'd906004072;
array2[8163]=30'd906004072;
array2[8164]=30'd906004072;
array2[8165]=30'd906004072;
array2[8166]=30'd906004072;
array2[8167]=30'd906004072;
array2[8168]=30'd906004072;
array2[8169]=30'd906004072;
array2[8170]=30'd906004072;
array2[8171]=30'd906004072;
array2[8172]=30'd906004072;
array2[8173]=30'd906004072;
array2[8174]=30'd906004072;
array2[8175]=30'd906004072;
array2[8176]=30'd906004072;
array2[8177]=30'd906004072;
array2[8178]=30'd906004072;
array2[8179]=30'd906004072;
array2[8180]=30'd906004072;
array2[8181]=30'd906004072;
array2[8182]=30'd906004072;
array2[8183]=30'd906004072;
array2[8184]=30'd906004072;
array2[8185]=30'd906004072;
array2[8186]=30'd906004072;
array2[8187]=30'd906004072;
array2[8188]=30'd906004072;
array2[8189]=30'd906004072;
array2[8190]=30'd906004072;
array2[8191]=30'd906004072;
array2[8192]=30'd906004072;
array2[8193]=30'd906004072;
array2[8194]=30'd906004072;
array2[8195]=30'd906004072;
array2[8196]=30'd906004072;
array2[8197]=30'd906004072;
array2[8198]=30'd906004072;
array2[8199]=30'd906004072;
array2[8200]=30'd906004072;
array2[8201]=30'd678604396;
array2[8202]=30'd538207812;
array2[8203]=30'd851505800;
array2[8204]=30'd851505800;
array2[8205]=30'd858839683;
array2[8206]=30'd851505800;
array2[8207]=30'd858839683;
array2[8208]=30'd858839683;
array2[8209]=30'd858839683;
array2[8210]=30'd865130113;
array2[8211]=30'd858839683;
array2[8212]=30'd865130113;
array2[8213]=30'd858839683;
array2[8214]=30'd858839683;
array2[8215]=30'd865130113;
array2[8216]=30'd858839683;
array2[8217]=30'd858839683;
array2[8218]=30'd858839683;
array2[8219]=30'd858839683;
array2[8220]=30'd858839683;
array2[8221]=30'd858839683;
array2[8222]=30'd851505800;
array2[8223]=30'd858839683;
array2[8224]=30'd858839683;
array2[8225]=30'd858839683;
array2[8226]=30'd858839683;
array2[8227]=30'd858839683;
array2[8228]=30'd851505800;
array2[8229]=30'd770812573;
array2[8230]=30'd828452495;
array2[8231]=30'd828452495;
array2[8232]=30'd506770009;
array2[8233]=30'd281508345;
array2[8234]=30'd764529268;
array2[8235]=30'd762499681;
array2[8236]=30'd281508345;
array2[8237]=30'd304706973;
array2[8238]=30'd312021416;
array2[8239]=30'd240774546;
array2[8240]=30'd227159434;
array2[8241]=30'd231362949;
array2[8242]=30'd231362949;
array2[8243]=30'd228216193;
array2[8244]=30'd229266819;
array2[8245]=30'd230317442;
array2[8246]=30'd229266819;
array2[8247]=30'd231364996;
array2[8248]=30'd231362949;
array2[8249]=30'd229266819;
array2[8250]=30'd229266819;
array2[8251]=30'd229266819;
array2[8252]=30'd229266819;
array2[8253]=30'd231362949;
array2[8254]=30'd229266819;
array2[8255]=30'd231362949;
array2[8256]=30'd790726247;
array2[8257]=30'd906004072;
array2[8258]=30'd906004072;
array2[8259]=30'd906004072;
array2[8260]=30'd736232864;
array2[8261]=30'd690121052;
array2[8262]=30'd690121052;
array2[8263]=30'd690121052;
array2[8264]=30'd690121052;
array2[8265]=30'd690121052;
array2[8266]=30'd690121052;
array2[8267]=30'd690121052;
array2[8268]=30'd690121052;
array2[8269]=30'd690121052;
array2[8270]=30'd690121052;
array2[8271]=30'd832648722;
array2[8272]=30'd906004072;
array2[8273]=30'd906004072;
array2[8274]=30'd906004072;
array2[8275]=30'd906004072;
array2[8276]=30'd906004072;
array2[8277]=30'd906004072;
array2[8278]=30'd906004072;
array2[8279]=30'd906004072;
array2[8280]=30'd906004072;
array2[8281]=30'd906004072;
array2[8282]=30'd906004072;
array2[8283]=30'd783393281;
array2[8284]=30'd690121052;
array2[8285]=30'd690121052;
array2[8286]=30'd690121052;
array2[8287]=30'd690121052;
array2[8288]=30'd690121052;
array2[8289]=30'd690121052;
array2[8290]=30'd690121052;
array2[8291]=30'd690121052;
array2[8292]=30'd690121052;
array2[8293]=30'd690121052;
array2[8294]=30'd783393281;
array2[8295]=30'd906004072;
array2[8296]=30'd823228019;
array2[8297]=30'd708987491;
array2[8298]=30'd538207812;
array2[8299]=30'd828452495;
array2[8300]=30'd858839683;
array2[8301]=30'd858839683;
array2[8302]=30'd851505800;
array2[8303]=30'd858839683;
array2[8304]=30'd851505800;
array2[8305]=30'd858839683;
array2[8306]=30'd858839683;
array2[8307]=30'd858839683;
array2[8308]=30'd865130113;
array2[8309]=30'd858839683;
array2[8310]=30'd858839683;
array2[8311]=30'd858839683;
array2[8312]=30'd858839683;
array2[8313]=30'd858839683;
array2[8314]=30'd858839683;
array2[8315]=30'd858839683;
array2[8316]=30'd858839683;
array2[8317]=30'd858839683;
array2[8318]=30'd865130113;
array2[8319]=30'd858839683;
array2[8320]=30'd858839683;
array2[8321]=30'd858839683;
array2[8322]=30'd858839683;
array2[8323]=30'd858839683;
array2[8324]=30'd828452495;
array2[8325]=30'd805398138;
array2[8326]=30'd828452495;
array2[8327]=30'd828452495;
array2[8328]=30'd506770009;
array2[8329]=30'd260631016;
array2[8330]=30'd790726247;
array2[8331]=30'd727851632;
array2[8332]=30'd281508345;
array2[8333]=30'd304706973;
array2[8334]=30'd271165847;
array2[8335]=30'd232392085;
array2[8336]=30'd227159434;
array2[8337]=30'd231362949;
array2[8338]=30'd231362949;
array2[8339]=30'd228216193;
array2[8340]=30'd229266819;
array2[8341]=30'd230317442;
array2[8342]=30'd231362949;
array2[8343]=30'd231362949;
array2[8344]=30'd229266819;
array2[8345]=30'd230317442;
array2[8346]=30'd231362949;
array2[8347]=30'd231364996;
array2[8348]=30'd229266819;
array2[8349]=30'd229266819;
array2[8350]=30'd228216193;
array2[8351]=30'd231362949;
array2[8352]=30'd639824186;
array2[8353]=30'd690121052;
array2[8354]=30'd690121052;
array2[8355]=30'd690121052;
array2[8356]=30'd637725975;
array2[8357]=30'd606284005;
array2[8358]=30'd606284005;
array2[8359]=30'd606284005;
array2[8360]=30'd606284005;
array2[8361]=30'd606284005;
array2[8362]=30'd606284005;
array2[8363]=30'd606284005;
array2[8364]=30'd606284005;
array2[8365]=30'd606284005;
array2[8366]=30'd611520752;
array2[8367]=30'd690121052;
array2[8368]=30'd690121052;
array2[8369]=30'd690121052;
array2[8370]=30'd690121052;
array2[8371]=30'd736232864;
array2[8372]=30'd690121052;
array2[8373]=30'd690121052;
array2[8374]=30'd690121052;
array2[8375]=30'd690121052;
array2[8376]=30'd690121052;
array2[8377]=30'd690121052;
array2[8378]=30'd736232864;
array2[8379]=30'd637725975;
array2[8380]=30'd611520752;
array2[8381]=30'd611520752;
array2[8382]=30'd611520752;
array2[8383]=30'd606284005;
array2[8384]=30'd606284005;
array2[8385]=30'd606284005;
array2[8386]=30'd606284005;
array2[8387]=30'd606284005;
array2[8388]=30'd606284005;
array2[8389]=30'd606284005;
array2[8390]=30'd639824186;
array2[8391]=30'd690121052;
array2[8392]=30'd690121052;
array2[8393]=30'd521469272;
array2[8394]=30'd506770009;
array2[8395]=30'd799112870;
array2[8396]=30'd828452495;
array2[8397]=30'd851505800;
array2[8398]=30'd858839683;
array2[8399]=30'd858839683;
array2[8400]=30'd858839683;
array2[8401]=30'd858839683;
array2[8402]=30'd858839683;
array2[8403]=30'd828452495;
array2[8404]=30'd770812573;
array2[8405]=30'd828452495;
array2[8406]=30'd828452495;
array2[8407]=30'd851505800;
array2[8408]=30'd851505800;
array2[8409]=30'd858839683;
array2[8410]=30'd851505800;
array2[8411]=30'd858839683;
array2[8412]=30'd851505800;
array2[8413]=30'd858839683;
array2[8414]=30'd858839683;
array2[8415]=30'd858839683;
array2[8416]=30'd858839683;
array2[8417]=30'd858839683;
array2[8418]=30'd858839683;
array2[8419]=30'd828452495;
array2[8420]=30'd732038833;
array2[8421]=30'd732038833;
array2[8422]=30'd799112870;
array2[8423]=30'd828452495;
array2[8424]=30'd566515308;
array2[8425]=30'd249001484;
array2[8426]=30'd764529268;
array2[8427]=30'd678602388;
array2[8428]=30'd281508345;
array2[8429]=30'd304706973;
array2[8430]=30'd257539480;
array2[8431]=30'd227159434;
array2[8432]=30'd227159434;
array2[8433]=30'd228216193;
array2[8434]=30'd230317442;
array2[8435]=30'd231364996;
array2[8436]=30'd231362949;
array2[8437]=30'd230317442;
array2[8438]=30'd229266819;
array2[8439]=30'd231362949;
array2[8440]=30'd229266819;
array2[8441]=30'd229266819;
array2[8442]=30'd229266819;
array2[8443]=30'd231359873;
array2[8444]=30'd231362949;
array2[8445]=30'd228216193;
array2[8446]=30'd227165569;
array2[8447]=30'd228216193;
array2[8448]=30'd582318295;
array2[8449]=30'd611520752;
array2[8450]=30'd611520752;
array2[8451]=30'd615715061;
array2[8452]=30'd611520752;
array2[8453]=30'd611520752;
array2[8454]=30'd611520752;
array2[8455]=30'd611520752;
array2[8456]=30'd611520752;
array2[8457]=30'd611520752;
array2[8458]=30'd611520752;
array2[8459]=30'd611520752;
array2[8460]=30'd611520752;
array2[8461]=30'd611520752;
array2[8462]=30'd611520752;
array2[8463]=30'd611520752;
array2[8464]=30'd606284005;
array2[8465]=30'd606284005;
array2[8466]=30'd611520752;
array2[8467]=30'd606284005;
array2[8468]=30'd606284005;
array2[8469]=30'd611520752;
array2[8470]=30'd611520752;
array2[8471]=30'd611520752;
array2[8472]=30'd611520752;
array2[8473]=30'd611520752;
array2[8474]=30'd611520752;
array2[8475]=30'd611520752;
array2[8476]=30'd611520752;
array2[8477]=30'd606284005;
array2[8478]=30'd611520752;
array2[8479]=30'd611520752;
array2[8480]=30'd611520752;
array2[8481]=30'd611520752;
array2[8482]=30'd611520752;
array2[8483]=30'd611520752;
array2[8484]=30'd611520752;
array2[8485]=30'd611520752;
array2[8486]=30'd606284005;
array2[8487]=30'd606284005;
array2[8488]=30'd595854564;
array2[8489]=30'd521469272;
array2[8490]=30'd449120871;
array2[8491]=30'd732038833;
array2[8492]=30'd828452495;
array2[8493]=30'd851505800;
array2[8494]=30'd851505800;
array2[8495]=30'd858839683;
array2[8496]=30'd858839683;
array2[8497]=30'd858839683;
array2[8498]=30'd858839683;
array2[8499]=30'd828452495;
array2[8500]=30'd678602388;
array2[8501]=30'd631447172;
array2[8502]=30'd727851632;
array2[8503]=30'd799112870;
array2[8504]=30'd828452495;
array2[8505]=30'd858839683;
array2[8506]=30'd851505800;
array2[8507]=30'd858839683;
array2[8508]=30'd858839683;
array2[8509]=30'd858839683;
array2[8510]=30'd858839683;
array2[8511]=30'd858839683;
array2[8512]=30'd858839683;
array2[8513]=30'd865130113;
array2[8514]=30'd851505800;
array2[8515]=30'd713202349;
array2[8516]=30'd409311115;
array2[8517]=30'd558174979;
array2[8518]=30'd646169309;
array2[8519]=30'd799112870;
array2[8520]=30'd560184961;
array2[8521]=30'd434416250;
array2[8522]=30'd764529268;
array2[8523]=30'd768729747;
array2[8524]=30'd506770009;
array2[8525]=30'd179916222;
array2[8526]=30'd212454818;
array2[8527]=30'd234504581;
array2[8528]=30'd231359873;
array2[8529]=30'd230317442;
array2[8530]=30'd231362949;
array2[8531]=30'd229266819;
array2[8532]=30'd231362949;
array2[8533]=30'd230317442;
array2[8534]=30'd231362949;
array2[8535]=30'd231362949;
array2[8536]=30'd231362949;
array2[8537]=30'd228216193;
array2[8538]=30'd229266819;
array2[8539]=30'd229266819;
array2[8540]=30'd230317442;
array2[8541]=30'd231362949;
array2[8542]=30'd227165569;
array2[8543]=30'd231362949;
array2[8544]=30'd582318295;
array2[8545]=30'd606284005;
array2[8546]=30'd611520752;
array2[8547]=30'd606284005;
array2[8548]=30'd586531028;
array2[8549]=30'd585627858;
array2[8550]=30'd585627858;
array2[8551]=30'd585627858;
array2[8552]=30'd585627858;
array2[8553]=30'd585627858;
array2[8554]=30'd585627858;
array2[8555]=30'd585627858;
array2[8556]=30'd585627858;
array2[8557]=30'd585627858;
array2[8558]=30'd585627858;
array2[8559]=30'd595854564;
array2[8560]=30'd611520752;
array2[8561]=30'd606284005;
array2[8562]=30'd606284005;
array2[8563]=30'd606284005;
array2[8564]=30'd611520752;
array2[8565]=30'd611520752;
array2[8566]=30'd606284005;
array2[8567]=30'd611520752;
array2[8568]=30'd611520752;
array2[8569]=30'd611520752;
array2[8570]=30'd606284005;
array2[8571]=30'd586531028;
array2[8572]=30'd585627858;
array2[8573]=30'd585627858;
array2[8574]=30'd585627858;
array2[8575]=30'd585627858;
array2[8576]=30'd585627858;
array2[8577]=30'd585627858;
array2[8578]=30'd585627858;
array2[8579]=30'd585627858;
array2[8580]=30'd585627858;
array2[8581]=30'd585627858;
array2[8582]=30'd586531028;
array2[8583]=30'd606284005;
array2[8584]=30'd595854564;
array2[8585]=30'd619916568;
array2[8586]=30'd521469272;
array2[8587]=30'd672348794;
array2[8588]=30'd770812573;
array2[8589]=30'd828452495;
array2[8590]=30'd851505800;
array2[8591]=30'd858839683;
array2[8592]=30'd858839683;
array2[8593]=30'd858839683;
array2[8594]=30'd865130113;
array2[8595]=30'd858839683;
array2[8596]=30'd828452495;
array2[8597]=30'd768729747;
array2[8598]=30'd631447172;
array2[8599]=30'd560184961;
array2[8600]=30'd711090860;
array2[8601]=30'd819020415;
array2[8602]=30'd851505800;
array2[8603]=30'd858839683;
array2[8604]=30'd851505800;
array2[8605]=30'd858839683;
array2[8606]=30'd858839683;
array2[8607]=30'd858839683;
array2[8608]=30'd858839683;
array2[8609]=30'd858839683;
array2[8610]=30'd711090860;
array2[8611]=30'd451191548;
array2[8612]=30'd451191548;
array2[8613]=30'd409311115;
array2[8614]=30'd558174979;
array2[8615]=30'd713179821;
array2[8616]=30'd805398138;
array2[8617]=30'd770816666;
array2[8618]=30'd828452495;
array2[8619]=30'd851505800;
array2[8620]=30'd770816666;
array2[8621]=30'd450208341;
array2[8622]=30'd207191473;
array2[8623]=30'd227165569;
array2[8624]=30'd231359873;
array2[8625]=30'd231362949;
array2[8626]=30'd229266819;
array2[8627]=30'd229266819;
array2[8628]=30'd231362949;
array2[8629]=30'd228216193;
array2[8630]=30'd231362949;
array2[8631]=30'd228216193;
array2[8632]=30'd228216193;
array2[8633]=30'd231359873;
array2[8634]=30'd231362949;
array2[8635]=30'd231362949;
array2[8636]=30'd229266819;
array2[8637]=30'd228216193;
array2[8638]=30'd228216193;
array2[8639]=30'd231362949;
array2[8640]=30'd561572038;
array2[8641]=30'd561572038;
array2[8642]=30'd561572038;
array2[8643]=30'd561572038;
array2[8644]=30'd514590904;
array2[8645]=30'd524037312;
array2[8646]=30'd518815920;
array2[8647]=30'd518815920;
array2[8648]=30'd518815920;
array2[8649]=30'd518815920;
array2[8650]=30'd518815920;
array2[8651]=30'd518815920;
array2[8652]=30'd518815920;
array2[8653]=30'd518815920;
array2[8654]=30'd524037312;
array2[8655]=30'd543866052;
array2[8656]=30'd561572038;
array2[8657]=30'd561572038;
array2[8658]=30'd561572038;
array2[8659]=30'd561572038;
array2[8660]=30'd561572038;
array2[8661]=30'd561572038;
array2[8662]=30'd561572038;
array2[8663]=30'd561572038;
array2[8664]=30'd561572038;
array2[8665]=30'd561572038;
array2[8666]=30'd561572038;
array2[8667]=30'd537610423;
array2[8668]=30'd524037312;
array2[8669]=30'd518815920;
array2[8670]=30'd518815920;
array2[8671]=30'd518815920;
array2[8672]=30'd518815920;
array2[8673]=30'd518815920;
array2[8674]=30'd518815920;
array2[8675]=30'd518815920;
array2[8676]=30'd518815920;
array2[8677]=30'd518815920;
array2[8678]=30'd537610423;
array2[8679]=30'd561572038;
array2[8680]=30'd561572038;
array2[8681]=30'd561572038;
array2[8682]=30'd452540782;
array2[8683]=30'd631447172;
array2[8684]=30'd732038833;
array2[8685]=30'd770812573;
array2[8686]=30'd828452495;
array2[8687]=30'd851505800;
array2[8688]=30'd851505800;
array2[8689]=30'd858839683;
array2[8690]=30'd858839683;
array2[8691]=30'd858839683;
array2[8692]=30'd865130113;
array2[8693]=30'd851505800;
array2[8694]=30'd828452495;
array2[8695]=30'd678602388;
array2[8696]=30'd560184961;
array2[8697]=30'd768729747;
array2[8698]=30'd828452495;
array2[8699]=30'd858839683;
array2[8700]=30'd858839683;
array2[8701]=30'd865130113;
array2[8702]=30'd858839683;
array2[8703]=30'd858839683;
array2[8704]=30'd858839683;
array2[8705]=30'd865130113;
array2[8706]=30'd601041592;
array2[8707]=30'd451191548;
array2[8708]=30'd451191548;
array2[8709]=30'd390446940;
array2[8710]=30'd409311115;
array2[8711]=30'd646169309;
array2[8712]=30'd858839683;
array2[8713]=30'd851505800;
array2[8714]=30'd819020415;
array2[8715]=30'd764529268;
array2[8716]=30'd713179821;
array2[8717]=30'd483727963;
array2[8718]=30'd193577377;
array2[8719]=30'd230307208;
array2[8720]=30'd228216193;
array2[8721]=30'd229266819;
array2[8722]=30'd228216193;
array2[8723]=30'd231359873;
array2[8724]=30'd231359873;
array2[8725]=30'd231362949;
array2[8726]=30'd231362949;
array2[8727]=30'd228216193;
array2[8728]=30'd231362949;
array2[8729]=30'd231362949;
array2[8730]=30'd231362949;
array2[8731]=30'd230317442;
array2[8732]=30'd230317442;
array2[8733]=30'd231362949;
array2[8734]=30'd228216193;
array2[8735]=30'd231364996;
array2[8736]=30'd496710898;
array2[8737]=30'd518815920;
array2[8738]=30'd518815920;
array2[8739]=30'd521966763;
array2[8740]=30'd521966763;
array2[8741]=30'd521966763;
array2[8742]=30'd521966763;
array2[8743]=30'd521966763;
array2[8744]=30'd521966763;
array2[8745]=30'd521966763;
array2[8746]=30'd521966763;
array2[8747]=30'd521966763;
array2[8748]=30'd521966763;
array2[8749]=30'd521966763;
array2[8750]=30'd521966763;
array2[8751]=30'd521966763;
array2[8752]=30'd518815920;
array2[8753]=30'd521966763;
array2[8754]=30'd521966763;
array2[8755]=30'd521966763;
array2[8756]=30'd521966763;
array2[8757]=30'd521966763;
array2[8758]=30'd521966763;
array2[8759]=30'd521966763;
array2[8760]=30'd518815920;
array2[8761]=30'd521966763;
array2[8762]=30'd518815920;
array2[8763]=30'd518815920;
array2[8764]=30'd521966763;
array2[8765]=30'd518815920;
array2[8766]=30'd521966763;
array2[8767]=30'd521966763;
array2[8768]=30'd521966763;
array2[8769]=30'd521966763;
array2[8770]=30'd521966763;
array2[8771]=30'd521966763;
array2[8772]=30'd521966763;
array2[8773]=30'd521966763;
array2[8774]=30'd521966763;
array2[8775]=30'd518815920;
array2[8776]=30'd518785242;
array2[8777]=30'd514590904;
array2[8778]=30'd498786593;
array2[8779]=30'd481587821;
array2[8780]=30'd678602388;
array2[8781]=30'd732038833;
array2[8782]=30'd770812573;
array2[8783]=30'd770812573;
array2[8784]=30'd828452495;
array2[8785]=30'd851505800;
array2[8786]=30'd858839683;
array2[8787]=30'd858839683;
array2[8788]=30'd858839683;
array2[8789]=30'd865130113;
array2[8790]=30'd858839683;
array2[8791]=30'd770812573;
array2[8792]=30'd560184961;
array2[8793]=30'd768729747;
array2[8794]=30'd828452495;
array2[8795]=30'd858839683;
array2[8796]=30'd858839683;
array2[8797]=30'd851505800;
array2[8798]=30'd858839683;
array2[8799]=30'd858839683;
array2[8800]=30'd858839683;
array2[8801]=30'd858839683;
array2[8802]=30'd770812573;
array2[8803]=30'd601041592;
array2[8804]=30'd451191548;
array2[8805]=30'd451191548;
array2[8806]=30'd601041592;
array2[8807]=30'd799112870;
array2[8808]=30'd819020415;
array2[8809]=30'd819020415;
array2[8810]=30'd764529268;
array2[8811]=30'd631447172;
array2[8812]=30'd483727963;
array2[8813]=30'd260631016;
array2[8814]=30'd228216193;
array2[8815]=30'd234504581;
array2[8816]=30'd229266819;
array2[8817]=30'd231362949;
array2[8818]=30'd230317442;
array2[8819]=30'd231362949;
array2[8820]=30'd229266819;
array2[8821]=30'd231362949;
array2[8822]=30'd230317442;
array2[8823]=30'd229266819;
array2[8824]=30'd229266819;
array2[8825]=30'd231362949;
array2[8826]=30'd229266819;
array2[8827]=30'd231362949;
array2[8828]=30'd231362949;
array2[8829]=30'd231362949;
array2[8830]=30'd231364996;
array2[8831]=30'd231362949;
array2[8832]=30'd496710898;
array2[8833]=30'd521966763;
array2[8834]=30'd521966763;
array2[8835]=30'd518815920;
array2[8836]=30'd515671261;
array2[8837]=30'd510427417;
array2[8838]=30'd510427417;
array2[8839]=30'd510427417;
array2[8840]=30'd510427417;
array2[8841]=30'd510427417;
array2[8842]=30'd510427417;
array2[8843]=30'd510427417;
array2[8844]=30'd510427417;
array2[8845]=30'd510427417;
array2[8846]=30'd510427417;
array2[8847]=30'd515671261;
array2[8848]=30'd521966763;
array2[8849]=30'd521966763;
array2[8850]=30'd521966763;
array2[8851]=30'd521966763;
array2[8852]=30'd521966763;
array2[8853]=30'd521966763;
array2[8854]=30'd521966763;
array2[8855]=30'd521966763;
array2[8856]=30'd521966763;
array2[8857]=30'd521966763;
array2[8858]=30'd521966763;
array2[8859]=30'd515671261;
array2[8860]=30'd510427417;
array2[8861]=30'd510427417;
array2[8862]=30'd510427417;
array2[8863]=30'd510427417;
array2[8864]=30'd510427417;
array2[8865]=30'd510427417;
array2[8866]=30'd510427417;
array2[8867]=30'd510427417;
array2[8868]=30'd510427417;
array2[8869]=30'd510427417;
array2[8870]=30'd515671261;
array2[8871]=30'd521966763;
array2[8872]=30'd524037312;
array2[8873]=30'd514590904;
array2[8874]=30'd537610423;
array2[8875]=30'd489282972;
array2[8876]=30'd506770009;
array2[8877]=30'd713202349;
array2[8878]=30'd732038833;
array2[8879]=30'd770812573;
array2[8880]=30'd770812573;
array2[8881]=30'd828452495;
array2[8882]=30'd851505800;
array2[8883]=30'd858839683;
array2[8884]=30'd858839683;
array2[8885]=30'd865130113;
array2[8886]=30'd828452495;
array2[8887]=30'd770812573;
array2[8888]=30'd560184961;
array2[8889]=30'd768729747;
array2[8890]=30'd828452495;
array2[8891]=30'd858839683;
array2[8892]=30'd858839683;
array2[8893]=30'd858839683;
array2[8894]=30'd858839683;
array2[8895]=30'd858839683;
array2[8896]=30'd858839683;
array2[8897]=30'd858839683;
array2[8898]=30'd858839683;
array2[8899]=30'd770816666;
array2[8900]=30'd646169309;
array2[8901]=30'd558174979;
array2[8902]=30'd768729747;
array2[8903]=30'd790726247;
array2[8904]=30'd790726247;
array2[8905]=30'd790726247;
array2[8906]=30'd764529268;
array2[8907]=30'd677571193;
array2[8908]=30'd506770009;
array2[8909]=30'd207191473;
array2[8910]=30'd231364996;
array2[8911]=30'd227165569;
array2[8912]=30'd231362949;
array2[8913]=30'd228216193;
array2[8914]=30'd229266819;
array2[8915]=30'd229266819;
array2[8916]=30'd231362949;
array2[8917]=30'd229266819;
array2[8918]=30'd229266819;
array2[8919]=30'd230317442;
array2[8920]=30'd231362949;
array2[8921]=30'd229266819;
array2[8922]=30'd231362949;
array2[8923]=30'd231362949;
array2[8924]=30'd229266819;
array2[8925]=30'd231362949;
array2[8926]=30'd231362949;
array2[8927]=30'd231364996;
array2[8928]=30'd387723742;
array2[8929]=30'd482131304;
array2[8930]=30'd482131304;
array2[8931]=30'd475838865;
array2[8932]=30'd473746934;
array2[8933]=30'd482138634;
array2[8934]=30'd475850257;
array2[8935]=30'd475850257;
array2[8936]=30'd475850257;
array2[8937]=30'd475850257;
array2[8938]=30'd475850257;
array2[8939]=30'd475850257;
array2[8940]=30'd475850257;
array2[8941]=30'd475850257;
array2[8942]=30'd482138634;
array2[8943]=30'd477946350;
array2[8944]=30'd482131304;
array2[8945]=30'd482131304;
array2[8946]=30'd482131304;
array2[8947]=30'd482131304;
array2[8948]=30'd482131304;
array2[8949]=30'd482131304;
array2[8950]=30'd482131304;
array2[8951]=30'd482131304;
array2[8952]=30'd482131304;
array2[8953]=30'd482131304;
array2[8954]=30'd482131304;
array2[8955]=30'd473746934;
array2[8956]=30'd482138634;
array2[8957]=30'd482138634;
array2[8958]=30'd482138634;
array2[8959]=30'd482138634;
array2[8960]=30'd480046615;
array2[8961]=30'd480046615;
array2[8962]=30'd480046615;
array2[8963]=30'd480046615;
array2[8964]=30'd480046615;
array2[8965]=30'd480046615;
array2[8966]=30'd477946350;
array2[8967]=30'd482131304;
array2[8968]=30'd475838865;
array2[8969]=30'd462205301;
array2[8970]=30'd528185854;
array2[8971]=30'd457992679;
array2[8972]=30'd425297329;
array2[8973]=30'd518272648;
array2[8974]=30'd713179821;
array2[8975]=30'd732038833;
array2[8976]=30'd770816666;
array2[8977]=30'd770812573;
array2[8978]=30'd799112870;
array2[8979]=30'd851505800;
array2[8980]=30'd851505800;
array2[8981]=30'd858839683;
array2[8982]=30'd770812573;
array2[8983]=30'd732038833;
array2[8984]=30'd560184961;
array2[8985]=30'd732038833;
array2[8986]=30'd819020415;
array2[8987]=30'd851505800;
array2[8988]=30'd828452495;
array2[8989]=30'd828452495;
array2[8990]=30'd851505800;
array2[8991]=30'd851505800;
array2[8992]=30'd828452495;
array2[8993]=30'd819020415;
array2[8994]=30'd828452495;
array2[8995]=30'd828452495;
array2[8996]=30'd819020415;
array2[8997]=30'd828452495;
array2[8998]=30'd828452495;
array2[8999]=30'd768729747;
array2[9000]=30'd764529268;
array2[9001]=30'd768729747;
array2[9002]=30'd678602388;
array2[9003]=30'd450208341;
array2[9004]=30'd195647926;
array2[9005]=30'd230307208;
array2[9006]=30'd231362949;
array2[9007]=30'd231359873;
array2[9008]=30'd231362949;
array2[9009]=30'd231362949;
array2[9010]=30'd231362949;
array2[9011]=30'd231362949;
array2[9012]=30'd229266819;
array2[9013]=30'd228216193;
array2[9014]=30'd231362949;
array2[9015]=30'd231362949;
array2[9016]=30'd229266819;
array2[9017]=30'd228216193;
array2[9018]=30'd229266819;
array2[9019]=30'd229266819;
array2[9020]=30'd231359873;
array2[9021]=30'd231364996;
array2[9022]=30'd227165569;
array2[9023]=30'd229266819;
array2[9024]=30'd387723742;
array2[9025]=30'd480046615;
array2[9026]=30'd480046615;
array2[9027]=30'd480046615;
array2[9028]=30'd480046615;
array2[9029]=30'd475850257;
array2[9030]=30'd475850257;
array2[9031]=30'd480046615;
array2[9032]=30'd480046615;
array2[9033]=30'd475850257;
array2[9034]=30'd480046615;
array2[9035]=30'd480046615;
array2[9036]=30'd475850257;
array2[9037]=30'd475850257;
array2[9038]=30'd475850257;
array2[9039]=30'd475850257;
array2[9040]=30'd475850257;
array2[9041]=30'd475850257;
array2[9042]=30'd475850257;
array2[9043]=30'd475850257;
array2[9044]=30'd482138634;
array2[9045]=30'd475850257;
array2[9046]=30'd482138634;
array2[9047]=30'd475850257;
array2[9048]=30'd482138634;
array2[9049]=30'd482138634;
array2[9050]=30'd475850257;
array2[9051]=30'd482138634;
array2[9052]=30'd475850257;
array2[9053]=30'd480046615;
array2[9054]=30'd475850257;
array2[9055]=30'd475850257;
array2[9056]=30'd480046615;
array2[9057]=30'd475850257;
array2[9058]=30'd480046615;
array2[9059]=30'd480046615;
array2[9060]=30'd480046615;
array2[9061]=30'd480046615;
array2[9062]=30'd480046615;
array2[9063]=30'd480046615;
array2[9064]=30'd480046615;
array2[9065]=30'd482138634;
array2[9066]=30'd509349393;
array2[9067]=30'd509349393;
array2[9068]=30'd509349393;
array2[9069]=30'd362496490;
array2[9070]=30'd449120871;
array2[9071]=30'd711090860;
array2[9072]=30'd770812573;
array2[9073]=30'd770812573;
array2[9074]=30'd770812573;
array2[9075]=30'd770812573;
array2[9076]=30'd770812573;
array2[9077]=30'd770812573;
array2[9078]=30'd732038833;
array2[9079]=30'd711090860;
array2[9080]=30'd678602388;
array2[9081]=30'd560184961;
array2[9082]=30'd518272648;
array2[9083]=30'd672348794;
array2[9084]=30'd805398138;
array2[9085]=30'd805398138;
array2[9086]=30'd805398138;
array2[9087]=30'd711090860;
array2[9088]=30'd732038833;
array2[9089]=30'd732038833;
array2[9090]=30'd770812573;
array2[9091]=30'd758240964;
array2[9092]=30'd770816666;
array2[9093]=30'd770812573;
array2[9094]=30'd770812573;
array2[9095]=30'd713179821;
array2[9096]=30'd678602388;
array2[9097]=30'd449120871;
array2[9098]=30'd347490866;
array2[9099]=30'd212454818;
array2[9100]=30'd231362949;
array2[9101]=30'd229266819;
array2[9102]=30'd229266819;
array2[9103]=30'd231362949;
array2[9104]=30'd231362949;
array2[9105]=30'd229266819;
array2[9106]=30'd231362949;
array2[9107]=30'd231362949;
array2[9108]=30'd231362949;
array2[9109]=30'd231362949;
array2[9110]=30'd229266819;
array2[9111]=30'd229266819;
array2[9112]=30'd230317442;
array2[9113]=30'd231362949;
array2[9114]=30'd231362949;
array2[9115]=30'd231362949;
array2[9116]=30'd231362949;
array2[9117]=30'd231362949;
array2[9118]=30'd231364996;
array2[9119]=30'd229266819;
array2[9120]=30'd439121402;
array2[9121]=30'd480046615;
array2[9122]=30'd480046615;
array2[9123]=30'd475850257;
array2[9124]=30'd439121402;
array2[9125]=30'd439121402;
array2[9126]=30'd387723742;
array2[9127]=30'd387723742;
array2[9128]=30'd387723742;
array2[9129]=30'd387723742;
array2[9130]=30'd387723742;
array2[9131]=30'd387723742;
array2[9132]=30'd387723742;
array2[9133]=30'd387723742;
array2[9134]=30'd387723742;
array2[9135]=30'd473746934;
array2[9136]=30'd475850257;
array2[9137]=30'd482138634;
array2[9138]=30'd482138634;
array2[9139]=30'd482138634;
array2[9140]=30'd482138634;
array2[9141]=30'd482138634;
array2[9142]=30'd482138634;
array2[9143]=30'd482138634;
array2[9144]=30'd482138634;
array2[9145]=30'd482138634;
array2[9146]=30'd482138634;
array2[9147]=30'd457992679;
array2[9148]=30'd387723742;
array2[9149]=30'd387723742;
array2[9150]=30'd387723742;
array2[9151]=30'd387723742;
array2[9152]=30'd387723742;
array2[9153]=30'd387723742;
array2[9154]=30'd387723742;
array2[9155]=30'd387723742;
array2[9156]=30'd439121402;
array2[9157]=30'd387723742;
array2[9158]=30'd457992679;
array2[9159]=30'd482138634;
array2[9160]=30'd475850257;
array2[9161]=30'd482138634;
array2[9162]=30'd482138634;
array2[9163]=30'd509349393;
array2[9164]=30'd509349393;
array2[9165]=30'd528185854;
array2[9166]=30'd362496490;
array2[9167]=30'd407216718;
array2[9168]=30'd407216718;
array2[9169]=30'd631447172;
array2[9170]=30'd770812573;
array2[9171]=30'd758240964;
array2[9172]=30'd732038833;
array2[9173]=30'd732038833;
array2[9174]=30'd732038833;
array2[9175]=30'd713179821;
array2[9176]=30'd560184961;
array2[9177]=30'd450208341;
array2[9178]=30'd407216718;
array2[9179]=30'd565444213;
array2[9180]=30'd790726247;
array2[9181]=30'd790726247;
array2[9182]=30'd711090860;
array2[9183]=30'd560184961;
array2[9184]=30'd678602388;
array2[9185]=30'd770816666;
array2[9186]=30'd770812573;
array2[9187]=30'd732038833;
array2[9188]=30'd732038833;
array2[9189]=30'd711090860;
array2[9190]=30'd518272648;
array2[9191]=30'd338018898;
array2[9192]=30'd319215128;
array2[9193]=30'd260631016;
array2[9194]=30'd228181405;
array2[9195]=30'd229266819;
array2[9196]=30'd231362949;
array2[9197]=30'd231364996;
array2[9198]=30'd231362949;
array2[9199]=30'd229266819;
array2[9200]=30'd231362949;
array2[9201]=30'd229266819;
array2[9202]=30'd229266819;
array2[9203]=30'd230317442;
array2[9204]=30'd229266819;
array2[9205]=30'd229266819;
array2[9206]=30'd231364996;
array2[9207]=30'd229266819;
array2[9208]=30'd229266819;
array2[9209]=30'd231362949;
array2[9210]=30'd231362949;
array2[9211]=30'd231364996;
array2[9212]=30'd231364996;
array2[9213]=30'd229266819;
array2[9214]=30'd228216193;
array2[9215]=30'd231364996;
array2[9216]=30'd362496490;
array2[9217]=30'd387723742;
array2[9218]=30'd387723742;
array2[9219]=30'd340509129;
array2[9220]=30'd302686639;
array2[9221]=30'd229270912;
array2[9222]=30'd234515845;
array2[9223]=30'd231364996;
array2[9224]=30'd228216193;
array2[9225]=30'd229270912;
array2[9226]=30'd232417668;
array2[9227]=30'd231362949;
array2[9228]=30'd229270912;
array2[9229]=30'd229270912;
array2[9230]=30'd232422779;
array2[9231]=30'd362496490;
array2[9232]=30'd387723742;
array2[9233]=30'd387723742;
array2[9234]=30'd387723742;
array2[9235]=30'd387723742;
array2[9236]=30'd387723742;
array2[9237]=30'd387723742;
array2[9238]=30'd387723742;
array2[9239]=30'd387723742;
array2[9240]=30'd387723742;
array2[9241]=30'd387723742;
array2[9242]=30'd340509129;
array2[9243]=30'd302686639;
array2[9244]=30'd234515845;
array2[9245]=30'd232434043;
array2[9246]=30'd232417668;
array2[9247]=30'd234515845;
array2[9248]=30'd234515845;
array2[9249]=30'd229270912;
array2[9250]=30'd229270912;
array2[9251]=30'd236604812;
array2[9252]=30'd228216193;
array2[9253]=30'd234515845;
array2[9254]=30'd307963313;
array2[9255]=30'd387723742;
array2[9256]=30'd387723742;
array2[9257]=30'd387723742;
array2[9258]=30'd387723742;
array2[9259]=30'd387723742;
array2[9260]=30'd387723742;
array2[9261]=30'd340509129;
array2[9262]=30'd362496490;
array2[9263]=30'd302686639;
array2[9264]=30'd267996623;
array2[9265]=30'd485780117;
array2[9266]=30'd713202349;
array2[9267]=30'd606320275;
array2[9268]=30'd383147560;
array2[9269]=30'd347490866;
array2[9270]=30'd347490866;
array2[9271]=30'd407216718;
array2[9272]=30'd606320275;
array2[9273]=30'd631447172;
array2[9274]=30'd672348794;
array2[9275]=30'd708987491;
array2[9276]=30'd790726247;
array2[9277]=30'd764529268;
array2[9278]=30'd566515308;
array2[9279]=30'd483727963;
array2[9280]=30'd481587821;
array2[9281]=30'd450208341;
array2[9282]=30'd383147560;
array2[9283]=30'd383147560;
array2[9284]=30'd319215128;
array2[9285]=30'd347490866;
array2[9286]=30'd260631016;
array2[9287]=30'd213516691;
array2[9288]=30'd220861839;
array2[9289]=30'd221916546;
array2[9290]=30'd228212100;
array2[9291]=30'd229266819;
array2[9292]=30'd229266819;
array2[9293]=30'd231362949;
array2[9294]=30'd231359873;
array2[9295]=30'd231362949;
array2[9296]=30'd231362949;
array2[9297]=30'd231362949;
array2[9298]=30'd231362949;
array2[9299]=30'd231359873;
array2[9300]=30'd231362949;
array2[9301]=30'd231364996;
array2[9302]=30'd230317442;
array2[9303]=30'd230317442;
array2[9304]=30'd231362949;
array2[9305]=30'd231362949;
array2[9306]=30'd231362949;
array2[9307]=30'd231362949;
array2[9308]=30'd229266819;
array2[9309]=30'd229266819;
array2[9310]=30'd231364996;
array2[9311]=30'd231364996;
array2[9312]=30'd193577377;
array2[9313]=30'd238691720;
array2[9314]=30'd228216193;
array2[9315]=30'd231362949;
array2[9316]=30'd229266819;
array2[9317]=30'd228216193;
array2[9318]=30'd231362949;
array2[9319]=30'd227165569;
array2[9320]=30'd231359873;
array2[9321]=30'd231362949;
array2[9322]=30'd231362949;
array2[9323]=30'd231359873;
array2[9324]=30'd229266819;
array2[9325]=30'd231359873;
array2[9326]=30'd229266819;
array2[9327]=30'd228216193;
array2[9328]=30'd231362949;
array2[9329]=30'd231362949;
array2[9330]=30'd227159434;
array2[9331]=30'd230307208;
array2[9332]=30'd227159434;
array2[9333]=30'd228216193;
array2[9334]=30'd229266819;
array2[9335]=30'd231362949;
array2[9336]=30'd229266819;
array2[9337]=30'd229266819;
array2[9338]=30'd231362949;
array2[9339]=30'd229266819;
array2[9340]=30'd231362949;
array2[9341]=30'd229266819;
array2[9342]=30'd231362949;
array2[9343]=30'd231362949;
array2[9344]=30'd228216193;
array2[9345]=30'd229266819;
array2[9346]=30'd231362949;
array2[9347]=30'd231362949;
array2[9348]=30'd231364996;
array2[9349]=30'd230317442;
array2[9350]=30'd231362949;
array2[9351]=30'd229266819;
array2[9352]=30'd227165569;
array2[9353]=30'd227165569;
array2[9354]=30'd231364996;
array2[9355]=30'd221916546;
array2[9356]=30'd228181405;
array2[9357]=30'd271165847;
array2[9358]=30'd280599950;
array2[9359]=30'd312021416;
array2[9360]=30'd260631016;
array2[9361]=30'd208120309;
array2[9362]=30'd249001484;
array2[9363]=30'd281508345;
array2[9364]=30'd295249323;
array2[9365]=30'd271165847;
array2[9366]=30'd227159434;
array2[9367]=30'd179916222;
array2[9368]=30'd560184961;
array2[9369]=30'd678602388;
array2[9370]=30'd727851632;
array2[9371]=30'd764529268;
array2[9372]=30'd790726247;
array2[9373]=30'd678604396;
array2[9374]=30'd506770009;
array2[9375]=30'd481587821;
array2[9376]=30'd407216718;
array2[9377]=30'd260631016;
array2[9378]=30'd295249323;
array2[9379]=30'd304706973;
array2[9380]=30'd257539480;
array2[9381]=30'd230307208;
array2[9382]=30'd230307208;
array2[9383]=30'd228216193;
array2[9384]=30'd228216193;
array2[9385]=30'd229266819;
array2[9386]=30'd229266819;
array2[9387]=30'd231362949;
array2[9388]=30'd231364996;
array2[9389]=30'd231362949;
array2[9390]=30'd231362949;
array2[9391]=30'd231362949;
array2[9392]=30'd230317442;
array2[9393]=30'd229266819;
array2[9394]=30'd230317442;
array2[9395]=30'd229266819;
array2[9396]=30'd229266819;
array2[9397]=30'd231362949;
array2[9398]=30'd229266819;
array2[9399]=30'd229266819;
array2[9400]=30'd229266819;
array2[9401]=30'd231362949;
array2[9402]=30'd229270912;
array2[9403]=30'd231362949;
array2[9404]=30'd229266819;
array2[9405]=30'd229266819;
array2[9406]=30'd231364996;
array2[9407]=30'd230317442;
array2[9408]=30'd193577377;
array2[9409]=30'd227165569;
array2[9410]=30'd228216193;
array2[9411]=30'd228216193;
array2[9412]=30'd230317442;
array2[9413]=30'd231364996;
array2[9414]=30'd229266819;
array2[9415]=30'd230317442;
array2[9416]=30'd229270912;
array2[9417]=30'd230317442;
array2[9418]=30'd231364996;
array2[9419]=30'd229270912;
array2[9420]=30'd229266819;
array2[9421]=30'd231362949;
array2[9422]=30'd229266819;
array2[9423]=30'd231359873;
array2[9424]=30'd231362949;
array2[9425]=30'd231362949;
array2[9426]=30'd231362949;
array2[9427]=30'd228216193;
array2[9428]=30'd229266819;
array2[9429]=30'd231362949;
array2[9430]=30'd231364996;
array2[9431]=30'd230317442;
array2[9432]=30'd230317442;
array2[9433]=30'd231362949;
array2[9434]=30'd229266819;
array2[9435]=30'd229266819;
array2[9436]=30'd231362949;
array2[9437]=30'd229266819;
array2[9438]=30'd231362949;
array2[9439]=30'd231362949;
array2[9440]=30'd231362949;
array2[9441]=30'd228216193;
array2[9442]=30'd231362949;
array2[9443]=30'd231362949;
array2[9444]=30'd231364996;
array2[9445]=30'd231362949;
array2[9446]=30'd229266819;
array2[9447]=30'd228216193;
array2[9448]=30'd231362949;
array2[9449]=30'd231362949;
array2[9450]=30'd234504581;
array2[9451]=30'd231362949;
array2[9452]=30'd228216193;
array2[9453]=30'd221916546;
array2[9454]=30'd280599950;
array2[9455]=30'd304706973;
array2[9456]=30'd304706973;
array2[9457]=30'd312021416;
array2[9458]=30'd312021416;
array2[9459]=30'd312021416;
array2[9460]=30'd304706973;
array2[9461]=30'd271165847;
array2[9462]=30'd227159434;
array2[9463]=30'd179916222;
array2[9464]=30'd606320275;
array2[9465]=30'd678602388;
array2[9466]=30'd764529268;
array2[9467]=30'd790726247;
array2[9468]=30'd764529268;
array2[9469]=30'd566515308;
array2[9470]=30'd518272648;
array2[9471]=30'd407216718;
array2[9472]=30'd195647926;
array2[9473]=30'd269069720;
array2[9474]=30'd280599950;
array2[9475]=30'd257539480;
array2[9476]=30'd227159434;
array2[9477]=30'd231364996;
array2[9478]=30'd231362949;
array2[9479]=30'd227165569;
array2[9480]=30'd229266819;
array2[9481]=30'd228216193;
array2[9482]=30'd231362949;
array2[9483]=30'd231359873;
array2[9484]=30'd229266819;
array2[9485]=30'd231362949;
array2[9486]=30'd229266819;
array2[9487]=30'd231359873;
array2[9488]=30'd231362949;
array2[9489]=30'd231362949;
array2[9490]=30'd229266819;
array2[9491]=30'd229266819;
array2[9492]=30'd231362949;
array2[9493]=30'd231362949;
array2[9494]=30'd231362949;
array2[9495]=30'd229266819;
array2[9496]=30'd231362949;
array2[9497]=30'd231362949;
array2[9498]=30'd231362949;
array2[9499]=30'd229270912;
array2[9500]=30'd231364996;
array2[9501]=30'd230317442;
array2[9502]=30'd231362949;
array2[9503]=30'd231364996;
array2[9504]=30'd193577377;
array2[9505]=30'd227165569;
array2[9506]=30'd228216193;
array2[9507]=30'd228216193;
array2[9508]=30'd230317442;
array2[9509]=30'd231364996;
array2[9510]=30'd228216193;
array2[9511]=30'd230317442;
array2[9512]=30'd232417668;
array2[9513]=30'd229266819;
array2[9514]=30'd231362949;
array2[9515]=30'd232417668;
array2[9516]=30'd229266819;
array2[9517]=30'd231362949;
array2[9518]=30'd228216193;
array2[9519]=30'd231359873;
array2[9520]=30'd228216193;
array2[9521]=30'd230317442;
array2[9522]=30'd231362949;
array2[9523]=30'd231362949;
array2[9524]=30'd231362949;
array2[9525]=30'd231362949;
array2[9526]=30'd230317442;
array2[9527]=30'd230317442;
array2[9528]=30'd230317442;
array2[9529]=30'd231362949;
array2[9530]=30'd230317442;
array2[9531]=30'd229266819;
array2[9532]=30'd231362949;
array2[9533]=30'd231362949;
array2[9534]=30'd228216193;
array2[9535]=30'd228216193;
array2[9536]=30'd231362949;
array2[9537]=30'd231362949;
array2[9538]=30'd231362949;
array2[9539]=30'd228216193;
array2[9540]=30'd227165569;
array2[9541]=30'd231362949;
array2[9542]=30'd231362949;
array2[9543]=30'd228216193;
array2[9544]=30'd231362949;
array2[9545]=30'd231364996;
array2[9546]=30'd231362949;
array2[9547]=30'd231362949;
array2[9548]=30'd229266819;
array2[9549]=30'd231362949;
array2[9550]=30'd220861839;
array2[9551]=30'd271165847;
array2[9552]=30'd280599950;
array2[9553]=30'd304706973;
array2[9554]=30'd312021416;
array2[9555]=30'd312021416;
array2[9556]=30'd271165847;
array2[9557]=30'd265928088;
array2[9558]=30'd234499470;
array2[9559]=30'd195647926;
array2[9560]=30'd606320275;
array2[9561]=30'd678602388;
array2[9562]=30'd764529268;
array2[9563]=30'd790726247;
array2[9564]=30'd677571193;
array2[9565]=30'd518272648;
array2[9566]=30'd485780117;
array2[9567]=30'd281508345;
array2[9568]=30'd232392085;
array2[9569]=30'd227159434;
array2[9570]=30'd265928088;
array2[9571]=30'd227159434;
array2[9572]=30'd234504581;
array2[9573]=30'd229266819;
array2[9574]=30'd229266819;
array2[9575]=30'd231362949;
array2[9576]=30'd229266819;
array2[9577]=30'd231362949;
array2[9578]=30'd231362949;
array2[9579]=30'd231362949;
array2[9580]=30'd229266819;
array2[9581]=30'd231362949;
array2[9582]=30'd229266819;
array2[9583]=30'd231362949;
array2[9584]=30'd231362949;
array2[9585]=30'd230317442;
array2[9586]=30'd229266819;
array2[9587]=30'd231362949;
array2[9588]=30'd231362949;
array2[9589]=30'd231364996;
array2[9590]=30'd231362949;
array2[9591]=30'd229266819;
array2[9592]=30'd231362949;
array2[9593]=30'd229270912;
array2[9594]=30'd231362949;
array2[9595]=30'd231364996;
array2[9596]=30'd231364996;
array2[9597]=30'd231362949;
array2[9598]=30'd231362949;
array2[9599]=30'd231362949;
array2[9600]=30'd193577377;
array2[9601]=30'd231359873;
array2[9602]=30'd227165569;
array2[9603]=30'd228216193;
array2[9604]=30'd230317442;
array2[9605]=30'd231362949;
array2[9606]=30'd229266819;
array2[9607]=30'd229270912;
array2[9608]=30'd234515845;
array2[9609]=30'd229266819;
array2[9610]=30'd231362949;
array2[9611]=30'd234515845;
array2[9612]=30'd230317442;
array2[9613]=30'd231362949;
array2[9614]=30'd229266819;
array2[9615]=30'd231359873;
array2[9616]=30'd229266819;
array2[9617]=30'd229266819;
array2[9618]=30'd231362949;
array2[9619]=30'd231362949;
array2[9620]=30'd234504581;
array2[9621]=30'd234504581;
array2[9622]=30'd229266819;
array2[9623]=30'd231364996;
array2[9624]=30'd231364996;
array2[9625]=30'd229266819;
array2[9626]=30'd231362949;
array2[9627]=30'd229266819;
array2[9628]=30'd231362949;
array2[9629]=30'd231362949;
array2[9630]=30'd229266819;
array2[9631]=30'd228216193;
array2[9632]=30'd229266819;
array2[9633]=30'd229266819;
array2[9634]=30'd231362949;
array2[9635]=30'd234504581;
array2[9636]=30'd227165569;
array2[9637]=30'd231362949;
array2[9638]=30'd231362949;
array2[9639]=30'd231362949;
array2[9640]=30'd228216193;
array2[9641]=30'd231362949;
array2[9642]=30'd230317442;
array2[9643]=30'd231362949;
array2[9644]=30'd234504581;
array2[9645]=30'd227165569;
array2[9646]=30'd238691720;
array2[9647]=30'd265928088;
array2[9648]=30'd271165847;
array2[9649]=30'd304706973;
array2[9650]=30'd280599950;
array2[9651]=30'd248105365;
array2[9652]=30'd221916546;
array2[9653]=30'd227165569;
array2[9654]=30'd238691720;
array2[9655]=30'd195647926;
array2[9656]=30'd606320275;
array2[9657]=30'd678602388;
array2[9658]=30'd764529268;
array2[9659]=30'd764529268;
array2[9660]=30'd565444213;
array2[9661]=30'd481587821;
array2[9662]=30'd338018898;
array2[9663]=30'd254365107;
array2[9664]=30'd221916546;
array2[9665]=30'd238691720;
array2[9666]=30'd238691720;
array2[9667]=30'd228216193;
array2[9668]=30'd231362949;
array2[9669]=30'd230317442;
array2[9670]=30'd229266819;
array2[9671]=30'd231362949;
array2[9672]=30'd231362949;
array2[9673]=30'd229266819;
array2[9674]=30'd231362949;
array2[9675]=30'd229266819;
array2[9676]=30'd229266819;
array2[9677]=30'd230317442;
array2[9678]=30'd229266819;
array2[9679]=30'd229266819;
array2[9680]=30'd231362949;
array2[9681]=30'd231362949;
array2[9682]=30'd229266819;
array2[9683]=30'd231362949;
array2[9684]=30'd231362949;
array2[9685]=30'd231364996;
array2[9686]=30'd231364996;
array2[9687]=30'd229266819;
array2[9688]=30'd228216193;
array2[9689]=30'd231362949;
array2[9690]=30'd230317442;
array2[9691]=30'd231362949;
array2[9692]=30'd231362949;
array2[9693]=30'd231364996;
array2[9694]=30'd231362949;
array2[9695]=30'd230317442;
array2[9696]=30'd193577377;
array2[9697]=30'd234504581;
array2[9698]=30'd227165569;
array2[9699]=30'd228216193;
array2[9700]=30'd230317442;
array2[9701]=30'd229266819;
array2[9702]=30'd229266819;
array2[9703]=30'd230317442;
array2[9704]=30'd229270912;
array2[9705]=30'd230317442;
array2[9706]=30'd231362949;
array2[9707]=30'd232417668;
array2[9708]=30'd230317442;
array2[9709]=30'd231362949;
array2[9710]=30'd231362949;
array2[9711]=30'd231362949;
array2[9712]=30'd229266819;
array2[9713]=30'd229266819;
array2[9714]=30'd231362949;
array2[9715]=30'd231362949;
array2[9716]=30'd231362949;
array2[9717]=30'd231362949;
array2[9718]=30'd229266819;
array2[9719]=30'd231362949;
array2[9720]=30'd231362949;
array2[9721]=30'd230317442;
array2[9722]=30'd229266819;
array2[9723]=30'd231362949;
array2[9724]=30'd231362949;
array2[9725]=30'd230317442;
array2[9726]=30'd230317442;
array2[9727]=30'd234504581;
array2[9728]=30'd230317442;
array2[9729]=30'd231362949;
array2[9730]=30'd229266819;
array2[9731]=30'd229266819;
array2[9732]=30'd231362949;
array2[9733]=30'd231362949;
array2[9734]=30'd231364996;
array2[9735]=30'd229266819;
array2[9736]=30'd229266819;
array2[9737]=30'd231362949;
array2[9738]=30'd231362949;
array2[9739]=30'd229266819;
array2[9740]=30'd231362949;
array2[9741]=30'd231364996;
array2[9742]=30'd234504581;
array2[9743]=30'd227159434;
array2[9744]=30'd257539480;
array2[9745]=30'd304706973;
array2[9746]=30'd295249323;
array2[9747]=30'd248105365;
array2[9748]=30'd221916546;
array2[9749]=30'd225072515;
array2[9750]=30'd227165569;
array2[9751]=30'd195647926;
array2[9752]=30'd518272648;
array2[9753]=30'd678602388;
array2[9754]=30'd764529268;
array2[9755]=30'd678604396;
array2[9756]=30'd518272648;
array2[9757]=30'd347490866;
array2[9758]=30'd212454818;
array2[9759]=30'd229266819;
array2[9760]=30'd229266819;
array2[9761]=30'd231362949;
array2[9762]=30'd229266819;
array2[9763]=30'd230317442;
array2[9764]=30'd234504581;
array2[9765]=30'd229266819;
array2[9766]=30'd229266819;
array2[9767]=30'd230317442;
array2[9768]=30'd229266819;
array2[9769]=30'd229266819;
array2[9770]=30'd231362949;
array2[9771]=30'd229266819;
array2[9772]=30'd229266819;
array2[9773]=30'd231362949;
array2[9774]=30'd231362949;
array2[9775]=30'd231364996;
array2[9776]=30'd229266819;
array2[9777]=30'd229266819;
array2[9778]=30'd229266819;
array2[9779]=30'd231362949;
array2[9780]=30'd230317442;
array2[9781]=30'd231362949;
array2[9782]=30'd231362949;
array2[9783]=30'd231362949;
array2[9784]=30'd231362949;
array2[9785]=30'd230317442;
array2[9786]=30'd231362949;
array2[9787]=30'd230317442;
array2[9788]=30'd231362949;
array2[9789]=30'd231362949;
array2[9790]=30'd230317442;
array2[9791]=30'd231362949;
array2[9792]=30'd193577377;
array2[9793]=30'd234504581;
array2[9794]=30'd227165569;
array2[9795]=30'd228216193;
array2[9796]=30'd230317442;
array2[9797]=30'd231362949;
array2[9798]=30'd229266819;
array2[9799]=30'd230317442;
array2[9800]=30'd232417668;
array2[9801]=30'd229266819;
array2[9802]=30'd231362949;
array2[9803]=30'd232417668;
array2[9804]=30'd229266819;
array2[9805]=30'd231362949;
array2[9806]=30'd229266819;
array2[9807]=30'd231359873;
array2[9808]=30'd229266819;
array2[9809]=30'd229266819;
array2[9810]=30'd234504581;
array2[9811]=30'd231362949;
array2[9812]=30'd231362949;
array2[9813]=30'd231362949;
array2[9814]=30'd230317442;
array2[9815]=30'd230317442;
array2[9816]=30'd231362949;
array2[9817]=30'd231362949;
array2[9818]=30'd229266819;
array2[9819]=30'd230317442;
array2[9820]=30'd231362949;
array2[9821]=30'd230317442;
array2[9822]=30'd230317442;
array2[9823]=30'd229266819;
array2[9824]=30'd229266819;
array2[9825]=30'd231362949;
array2[9826]=30'd231362949;
array2[9827]=30'd229266819;
array2[9828]=30'd231362949;
array2[9829]=30'd231362949;
array2[9830]=30'd231362949;
array2[9831]=30'd230317442;
array2[9832]=30'd231362949;
array2[9833]=30'd231362949;
array2[9834]=30'd231362949;
array2[9835]=30'd230317442;
array2[9836]=30'd231362949;
array2[9837]=30'd234504581;
array2[9838]=30'd231362949;
array2[9839]=30'd234504581;
array2[9840]=30'd227165569;
array2[9841]=30'd248105365;
array2[9842]=30'd280599950;
array2[9843]=30'd271165847;
array2[9844]=30'd257539480;
array2[9845]=30'd227159434;
array2[9846]=30'd227165569;
array2[9847]=30'd221916546;
array2[9848]=30'd319215128;
array2[9849]=30'd560184961;
array2[9850]=30'd678602388;
array2[9851]=30'd565444213;
array2[9852]=30'd450208341;
array2[9853]=30'd265736724;
array2[9854]=30'd220861839;
array2[9855]=30'd228216193;
array2[9856]=30'd229266819;
array2[9857]=30'd231364996;
array2[9858]=30'd228216193;
array2[9859]=30'd229266819;
array2[9860]=30'd231362949;
array2[9861]=30'd229266819;
array2[9862]=30'd230317442;
array2[9863]=30'd230317442;
array2[9864]=30'd229266819;
array2[9865]=30'd229266819;
array2[9866]=30'd231364996;
array2[9867]=30'd229266819;
array2[9868]=30'd229266819;
array2[9869]=30'd231362949;
array2[9870]=30'd228216193;
array2[9871]=30'd231364996;
array2[9872]=30'd229266819;
array2[9873]=30'd229266819;
array2[9874]=30'd228216193;
array2[9875]=30'd228216193;
array2[9876]=30'd230317442;
array2[9877]=30'd231362949;
array2[9878]=30'd231362949;
array2[9879]=30'd231362949;
array2[9880]=30'd231362949;
array2[9881]=30'd230317442;
array2[9882]=30'd231362949;
array2[9883]=30'd231362949;
array2[9884]=30'd227165569;
array2[9885]=30'd231362949;
array2[9886]=30'd230317442;
array2[9887]=30'd229266819;
array2[9888]=30'd193577377;
array2[9889]=30'd234504581;
array2[9890]=30'd227165569;
array2[9891]=30'd228216193;
array2[9892]=30'd229266819;
array2[9893]=30'd229266819;
array2[9894]=30'd229266819;
array2[9895]=30'd230317442;
array2[9896]=30'd229270912;
array2[9897]=30'd229266819;
array2[9898]=30'd231362949;
array2[9899]=30'd229270912;
array2[9900]=30'd231362949;
array2[9901]=30'd231359873;
array2[9902]=30'd229266819;
array2[9903]=30'd231359873;
array2[9904]=30'd229266819;
array2[9905]=30'd228216193;
array2[9906]=30'd231362949;
array2[9907]=30'd231362949;
array2[9908]=30'd231362949;
array2[9909]=30'd231362949;
array2[9910]=30'd230317442;
array2[9911]=30'd231362949;
array2[9912]=30'd229266819;
array2[9913]=30'd231364996;
array2[9914]=30'd228216193;
array2[9915]=30'd231362949;
array2[9916]=30'd231362949;
array2[9917]=30'd231364996;
array2[9918]=30'd229266819;
array2[9919]=30'd228216193;
array2[9920]=30'd231362949;
array2[9921]=30'd231362949;
array2[9922]=30'd231362949;
array2[9923]=30'd231364996;
array2[9924]=30'd231362949;
array2[9925]=30'd231362949;
array2[9926]=30'd228216193;
array2[9927]=30'd231362949;
array2[9928]=30'd234504581;
array2[9929]=30'd231362949;
array2[9930]=30'd231362949;
array2[9931]=30'd229266819;
array2[9932]=30'd229266819;
array2[9933]=30'd231359873;
array2[9934]=30'd231362949;
array2[9935]=30'd231362949;
array2[9936]=30'd231362949;
array2[9937]=30'd231362949;
array2[9938]=30'd238691720;
array2[9939]=30'd221916546;
array2[9940]=30'd227159434;
array2[9941]=30'd227159434;
array2[9942]=30'd227165569;
array2[9943]=30'd231362949;
array2[9944]=30'd381167075;
array2[9945]=30'd281508345;
array2[9946]=30'd401997362;
array2[9947]=30'd319215128;
array2[9948]=30'd319215128;
array2[9949]=30'd190356956;
array2[9950]=30'd213516691;
array2[9951]=30'd229266819;
array2[9952]=30'd231364996;
array2[9953]=30'd231364996;
array2[9954]=30'd228216193;
array2[9955]=30'd229266819;
array2[9956]=30'd231362949;
array2[9957]=30'd231362949;
array2[9958]=30'd230317442;
array2[9959]=30'd231362949;
array2[9960]=30'd231362949;
array2[9961]=30'd231359873;
array2[9962]=30'd228216193;
array2[9963]=30'd231362949;
array2[9964]=30'd234504581;
array2[9965]=30'd231362949;
array2[9966]=30'd227165569;
array2[9967]=30'd229266819;
array2[9968]=30'd230317442;
array2[9969]=30'd231364996;
array2[9970]=30'd231362949;
array2[9971]=30'd227165569;
array2[9972]=30'd229266819;
array2[9973]=30'd228216193;
array2[9974]=30'd231362949;
array2[9975]=30'd228216193;
array2[9976]=30'd229266819;
array2[9977]=30'd229266819;
array2[9978]=30'd231359873;
array2[9979]=30'd231362949;
array2[9980]=30'd230307208;
array2[9981]=30'd227165569;
array2[9982]=30'd231362949;
array2[9983]=30'd229266819;
array2[9984]=30'd193577377;
array2[9985]=30'd234504581;
array2[9986]=30'd227165569;
array2[9987]=30'd228216193;
array2[9988]=30'd230317442;
array2[9989]=30'd231362949;
array2[9990]=30'd229266819;
array2[9991]=30'd229270912;
array2[9992]=30'd232417668;
array2[9993]=30'd229266819;
array2[9994]=30'd231362949;
array2[9995]=30'd234515845;
array2[9996]=30'd229266819;
array2[9997]=30'd231362949;
array2[9998]=30'd256519562;
array2[9999]=30'd231364996;
array2[10000]=30'd231362949;
array2[10001]=30'd231362949;
array2[10002]=30'd228212100;
array2[10003]=30'd231362949;
array2[10004]=30'd228216193;
array2[10005]=30'd231362949;
array2[10006]=30'd230317442;
array2[10007]=30'd231362949;
array2[10008]=30'd231362949;
array2[10009]=30'd231362949;
array2[10010]=30'd231362949;
array2[10011]=30'd231362949;
array2[10012]=30'd231362949;
array2[10013]=30'd231362949;
array2[10014]=30'd229266819;
array2[10015]=30'd228216193;
array2[10016]=30'd231362949;
array2[10017]=30'd231362949;
array2[10018]=30'd231362949;
array2[10019]=30'd231362949;
array2[10020]=30'd229266819;
array2[10021]=30'd256519562;
array2[10022]=30'd236604812;
array2[10023]=30'd231364996;
array2[10024]=30'd231362949;
array2[10025]=30'd229266819;
array2[10026]=30'd231362949;
array2[10027]=30'd231364996;
array2[10028]=30'd231364996;
array2[10029]=30'd229266819;
array2[10030]=30'd230317442;
array2[10031]=30'd231362949;
array2[10032]=30'd301610387;
array2[10033]=30'd272255371;
array2[10034]=30'd229266819;
array2[10035]=30'd229266819;
array2[10036]=30'd231362949;
array2[10037]=30'd229266819;
array2[10038]=30'd229266819;
array2[10039]=30'd231362949;
array2[10040]=30'd238691720;
array2[10041]=30'd227159434;
array2[10042]=30'd238691720;
array2[10043]=30'd227159434;
array2[10044]=30'd238691720;
array2[10045]=30'd230307208;
array2[10046]=30'd225072515;
array2[10047]=30'd229266819;
array2[10048]=30'd231362949;
array2[10049]=30'd231364996;
array2[10050]=30'd231362949;
array2[10051]=30'd230317442;
array2[10052]=30'd231362949;
array2[10053]=30'd230317442;
array2[10054]=30'd231362949;
array2[10055]=30'd231362949;
array2[10056]=30'd229266819;
array2[10057]=30'd231362949;
array2[10058]=30'd230317442;
array2[10059]=30'd231362949;
array2[10060]=30'd231364996;
array2[10061]=30'd231362949;
array2[10062]=30'd229266819;
array2[10063]=30'd231362949;
array2[10064]=30'd229266819;
array2[10065]=30'd229266819;
array2[10066]=30'd231362949;
array2[10067]=30'd229266819;
array2[10068]=30'd229266819;
array2[10069]=30'd231362949;
array2[10070]=30'd229266819;
array2[10071]=30'd231362949;
array2[10072]=30'd231362949;
array2[10073]=30'd231362949;
array2[10074]=30'd230317442;
array2[10075]=30'd231362949;
array2[10076]=30'd231362949;
array2[10077]=30'd228216193;
array2[10078]=30'd230317442;
array2[10079]=30'd230317442;
array2[10080]=30'd193577377;
array2[10081]=30'd234504581;
array2[10082]=30'd227165569;
array2[10083]=30'd228216193;
array2[10084]=30'd230317442;
array2[10085]=30'd229266819;
array2[10086]=30'd229266819;
array2[10087]=30'd230317442;
array2[10088]=30'd229270912;
array2[10089]=30'd229266819;
array2[10090]=30'd231362949;
array2[10091]=30'd229270912;
array2[10092]=30'd230317442;
array2[10093]=30'd272255371;
array2[10094]=30'd472496545;
array2[10095]=30'd272255371;
array2[10096]=30'd225072515;
array2[10097]=30'd231362949;
array2[10098]=30'd228216193;
array2[10099]=30'd228216193;
array2[10100]=30'd228216193;
array2[10101]=30'd231362949;
array2[10102]=30'd229266819;
array2[10103]=30'd231362949;
array2[10104]=30'd231362949;
array2[10105]=30'd231362949;
array2[10106]=30'd230317442;
array2[10107]=30'd231362949;
array2[10108]=30'd231362949;
array2[10109]=30'd229266819;
array2[10110]=30'd230317442;
array2[10111]=30'd229266819;
array2[10112]=30'd230317442;
array2[10113]=30'd231362949;
array2[10114]=30'd231364996;
array2[10115]=30'd231362949;
array2[10116]=30'd231362949;
array2[10117]=30'd405404052;
array2[10118]=30'd338288022;
array2[10119]=30'd228212100;
array2[10120]=30'd229270912;
array2[10121]=30'd228216193;
array2[10122]=30'd231364996;
array2[10123]=30'd230317442;
array2[10124]=30'd231362949;
array2[10125]=30'd231364996;
array2[10126]=30'd230317442;
array2[10127]=30'd256519562;
array2[10128]=30'd664345022;
array2[10129]=30'd553231776;
array2[10130]=30'd228212100;
array2[10131]=30'd229266819;
array2[10132]=30'd231362949;
array2[10133]=30'd228216193;
array2[10134]=30'd231359873;
array2[10135]=30'd231362949;
array2[10136]=30'd230317442;
array2[10137]=30'd230317442;
array2[10138]=30'd231362949;
array2[10139]=30'd229266819;
array2[10140]=30'd229266819;
array2[10141]=30'd231362949;
array2[10142]=30'd231362949;
array2[10143]=30'd229266819;
array2[10144]=30'd229266819;
array2[10145]=30'd229266819;
array2[10146]=30'd229266819;
array2[10147]=30'd231362949;
array2[10148]=30'd231362949;
array2[10149]=30'd228216193;
array2[10150]=30'd229266819;
array2[10151]=30'd231362949;
array2[10152]=30'd231362949;
array2[10153]=30'd231364996;
array2[10154]=30'd229266819;
array2[10155]=30'd229266819;
array2[10156]=30'd231362949;
array2[10157]=30'd231362949;
array2[10158]=30'd227165569;
array2[10159]=30'd234504581;
array2[10160]=30'd231364996;
array2[10161]=30'd231362949;
array2[10162]=30'd231364996;
array2[10163]=30'd229266819;
array2[10164]=30'd231362949;
array2[10165]=30'd231362949;
array2[10166]=30'd231362949;
array2[10167]=30'd231362949;
array2[10168]=30'd231362949;
array2[10169]=30'd230317442;
array2[10170]=30'd229266819;
array2[10171]=30'd228216193;
array2[10172]=30'd231362949;
array2[10173]=30'd229266819;
array2[10174]=30'd229266819;
array2[10175]=30'd231362949;
array2[10176]=30'd193577377;
array2[10177]=30'd234504581;
array2[10178]=30'd227165569;
array2[10179]=30'd228216193;
array2[10180]=30'd230317442;
array2[10181]=30'd229266819;
array2[10182]=30'd229266819;
array2[10183]=30'd230317442;
array2[10184]=30'd229270912;
array2[10185]=30'd229266819;
array2[10186]=30'd231362949;
array2[10187]=30'd405404052;
array2[10188]=30'd338288022;
array2[10189]=30'd231362949;
array2[10190]=30'd272255371;
array2[10191]=30'd234504581;
array2[10192]=30'd272255371;
array2[10193]=30'd405404052;
array2[10194]=30'd231362949;
array2[10195]=30'd231362949;
array2[10196]=30'd231362949;
array2[10197]=30'd231362949;
array2[10198]=30'd231359873;
array2[10199]=30'd231359873;
array2[10200]=30'd231362949;
array2[10201]=30'd231362949;
array2[10202]=30'd228216193;
array2[10203]=30'd228216193;
array2[10204]=30'd231362949;
array2[10205]=30'd231362949;
array2[10206]=30'd231362949;
array2[10207]=30'd230317442;
array2[10208]=30'd230317442;
array2[10209]=30'd231362949;
array2[10210]=30'd377085336;
array2[10211]=30'd377085336;
array2[10212]=30'd230307208;
array2[10213]=30'd262793620;
array2[10214]=30'd231362949;
array2[10215]=30'd229266819;
array2[10216]=30'd428475791;
array2[10217]=30'd272255371;
array2[10218]=30'd234504581;
array2[10219]=30'd231362949;
array2[10220]=30'd231364996;
array2[10221]=30'd231364996;
array2[10222]=30'd231362949;
array2[10223]=30'd234504581;
array2[10224]=30'd272255371;
array2[10225]=30'd256519562;
array2[10226]=30'd228216193;
array2[10227]=30'd231362949;
array2[10228]=30'd228216193;
array2[10229]=30'd231362949;
array2[10230]=30'd231359873;
array2[10231]=30'd231362949;
array2[10232]=30'd231362949;
array2[10233]=30'd229266819;
array2[10234]=30'd228216193;
array2[10235]=30'd231362949;
array2[10236]=30'd231364996;
array2[10237]=30'd231362949;
array2[10238]=30'd229266819;
array2[10239]=30'd229266819;
array2[10240]=30'd231364996;
array2[10241]=30'd229266819;
array2[10242]=30'd231364996;
array2[10243]=30'd231362949;
array2[10244]=30'd231362949;
array2[10245]=30'd229266819;
array2[10246]=30'd229266819;
array2[10247]=30'd231362949;
array2[10248]=30'd234504581;
array2[10249]=30'd231362949;
array2[10250]=30'd228216193;
array2[10251]=30'd228216193;
array2[10252]=30'd231362949;
array2[10253]=30'd231362949;
array2[10254]=30'd227165569;
array2[10255]=30'd229266819;
array2[10256]=30'd229266819;
array2[10257]=30'd230317442;
array2[10258]=30'd231362949;
array2[10259]=30'd231362949;
array2[10260]=30'd231362949;
array2[10261]=30'd231362949;
array2[10262]=30'd231362949;
array2[10263]=30'd229266819;
array2[10264]=30'd231359873;
array2[10265]=30'd231364996;
array2[10266]=30'd230317442;
array2[10267]=30'd229266819;
array2[10268]=30'd230317442;
array2[10269]=30'd231362949;
array2[10270]=30'd231359873;
array2[10271]=30'd231362949;
array2[10272]=30'd193577377;
array2[10273]=30'd227165569;
array2[10274]=30'd227165569;
array2[10275]=30'd231362949;
array2[10276]=30'd229266819;
array2[10277]=30'd230317442;
array2[10278]=30'd231362949;
array2[10279]=30'd228216193;
array2[10280]=30'd229266819;
array2[10281]=30'd229266819;
array2[10282]=30'd229270912;
array2[10283]=30'd234504581;
array2[10284]=30'd231362949;
array2[10285]=30'd229270912;
array2[10286]=30'd230317442;
array2[10287]=30'd231362949;
array2[10288]=30'd231362949;
array2[10289]=30'd229270912;
array2[10290]=30'd229270912;
array2[10291]=30'd227165569;
array2[10292]=30'd231364996;
array2[10293]=30'd238691720;
array2[10294]=30'd234504581;
array2[10295]=30'd229266819;
array2[10296]=30'd231362949;
array2[10297]=30'd231362949;
array2[10298]=30'd228216193;
array2[10299]=30'd231362949;
array2[10300]=30'd231359873;
array2[10301]=30'd231362949;
array2[10302]=30'd228216193;
array2[10303]=30'd230317442;
array2[10304]=30'd229266819;
array2[10305]=30'd256519562;
array2[10306]=30'd236604812;
array2[10307]=30'd234504581;
array2[10308]=30'd231362949;
array2[10309]=30'd231362949;
array2[10310]=30'd229270912;
array2[10311]=30'd228216193;
array2[10312]=30'd236604812;
array2[10313]=30'd229270912;
array2[10314]=30'd227165569;
array2[10315]=30'd231362949;
array2[10316]=30'd234504581;
array2[10317]=30'd236604812;
array2[10318]=30'd231362949;
array2[10319]=30'd231362949;
array2[10320]=30'd231362949;
array2[10321]=30'd229270912;
array2[10322]=30'd231362949;
array2[10323]=30'd231362949;
array2[10324]=30'd231362949;
array2[10325]=30'd234499470;
array2[10326]=30'd228216193;
array2[10327]=30'd231359873;
array2[10328]=30'd231359873;
array2[10329]=30'd231362949;
array2[10330]=30'd230317442;
array2[10331]=30'd230317442;
array2[10332]=30'd231362949;
array2[10333]=30'd229266819;
array2[10334]=30'd229266819;
array2[10335]=30'd231362949;
array2[10336]=30'd231362949;
array2[10337]=30'd229266819;
array2[10338]=30'd228216193;
array2[10339]=30'd228216193;
array2[10340]=30'd229266819;
array2[10341]=30'd231359873;
array2[10342]=30'd234504581;
array2[10343]=30'd227165569;
array2[10344]=30'd227165569;
array2[10345]=30'd231362949;
array2[10346]=30'd234504581;
array2[10347]=30'd228216193;
array2[10348]=30'd228216193;
array2[10349]=30'd229266819;
array2[10350]=30'd231362949;
array2[10351]=30'd228216193;
array2[10352]=30'd227165569;
array2[10353]=30'd230307208;
array2[10354]=30'd231362949;
array2[10355]=30'd229266819;
array2[10356]=30'd231364996;
array2[10357]=30'd231362949;
array2[10358]=30'd231364996;
array2[10359]=30'd230317442;
array2[10360]=30'd231362949;
array2[10361]=30'd231362949;
array2[10362]=30'd229266819;
array2[10363]=30'd229266819;
array2[10364]=30'd229266819;
array2[10365]=30'd229266819;
array2[10366]=30'd231362949;
array2[10367]=30'd231362949;
array2[10368]=30'd212454818;
array2[10369]=30'd234504581;
array2[10370]=30'd231362949;
array2[10371]=30'd230317442;
array2[10372]=30'd229266819;
array2[10373]=30'd231362949;
array2[10374]=30'd231362949;
array2[10375]=30'd231362949;
array2[10376]=30'd231362949;
array2[10377]=30'd231362949;
array2[10378]=30'd231362949;
array2[10379]=30'd231359873;
array2[10380]=30'd229270912;
array2[10381]=30'd231362949;
array2[10382]=30'd228216193;
array2[10383]=30'd231364996;
array2[10384]=30'd229266819;
array2[10385]=30'd231362949;
array2[10386]=30'd231362949;
array2[10387]=30'd231362949;
array2[10388]=30'd231362949;
array2[10389]=30'd231362949;
array2[10390]=30'd231364996;
array2[10391]=30'd229266819;
array2[10392]=30'd229270912;
array2[10393]=30'd231362949;
array2[10394]=30'd231362949;
array2[10395]=30'd231362949;
array2[10396]=30'd230317442;
array2[10397]=30'd229266819;
array2[10398]=30'd229266819;
array2[10399]=30'd231362949;
array2[10400]=30'd234504581;
array2[10401]=30'd231362949;
array2[10402]=30'd231362949;
array2[10403]=30'd231362949;
array2[10404]=30'd231362949;
array2[10405]=30'd232417668;
array2[10406]=30'd231364996;
array2[10407]=30'd234504581;
array2[10408]=30'd231364996;
array2[10409]=30'd230317442;
array2[10410]=30'd229266819;
array2[10411]=30'd231362949;
array2[10412]=30'd231359873;
array2[10413]=30'd228216193;
array2[10414]=30'd231362949;
array2[10415]=30'd231362949;
array2[10416]=30'd231362949;
array2[10417]=30'd231362949;
array2[10418]=30'd229270912;
array2[10419]=30'd229266819;
array2[10420]=30'd229266819;
array2[10421]=30'd231362949;
array2[10422]=30'd228216193;
array2[10423]=30'd231362949;
array2[10424]=30'd229266819;
array2[10425]=30'd231362949;
array2[10426]=30'd229266819;
array2[10427]=30'd231364996;
array2[10428]=30'd231362949;
array2[10429]=30'd234504581;
array2[10430]=30'd231362949;
array2[10431]=30'd231359873;
array2[10432]=30'd229266819;
array2[10433]=30'd230317442;
array2[10434]=30'd231362949;
array2[10435]=30'd231362949;
array2[10436]=30'd228216193;
array2[10437]=30'd229266819;
array2[10438]=30'd231362949;
array2[10439]=30'd231362949;
array2[10440]=30'd231362949;
array2[10441]=30'd231362949;
array2[10442]=30'd231362949;
array2[10443]=30'd231362949;
array2[10444]=30'd229266819;
array2[10445]=30'd231364996;
array2[10446]=30'd229270912;
array2[10447]=30'd231362949;
array2[10448]=30'd377085336;
array2[10449]=30'd272255371;
array2[10450]=30'd338288022;
array2[10451]=30'd664345022;
array2[10452]=30'd338288022;
array2[10453]=30'd256519562;
array2[10454]=30'd377085336;
array2[10455]=30'd231362949;
array2[10456]=30'd230317442;
array2[10457]=30'd230317442;
array2[10458]=30'd229266819;
array2[10459]=30'd228216193;
array2[10460]=30'd231362949;
array2[10461]=30'd231362949;
array2[10462]=30'd231362949;
array2[10463]=30'd231362949;
array2[10464]=30'd193577377;
array2[10465]=30'd227165569;
array2[10466]=30'd228216193;
array2[10467]=30'd227165569;
array2[10468]=30'd231362949;
array2[10469]=30'd231362949;
array2[10470]=30'd229266819;
array2[10471]=30'd229266819;
array2[10472]=30'd228216193;
array2[10473]=30'd231364996;
array2[10474]=30'd229266819;
array2[10475]=30'd229266819;
array2[10476]=30'd229266819;
array2[10477]=30'd229266819;
array2[10478]=30'd231362949;
array2[10479]=30'd231362949;
array2[10480]=30'd229266819;
array2[10481]=30'd231362949;
array2[10482]=30'd230317442;
array2[10483]=30'd230317442;
array2[10484]=30'd229266819;
array2[10485]=30'd229266819;
array2[10486]=30'd231362949;
array2[10487]=30'd231362949;
array2[10488]=30'd231362949;
array2[10489]=30'd231362949;
array2[10490]=30'd231362949;
array2[10491]=30'd229266819;
array2[10492]=30'd231362949;
array2[10493]=30'd231362949;
array2[10494]=30'd231362949;
array2[10495]=30'd228216193;
array2[10496]=30'd231362949;
array2[10497]=30'd229266819;
array2[10498]=30'd231362949;
array2[10499]=30'd231364996;
array2[10500]=30'd234504581;
array2[10501]=30'd231362949;
array2[10502]=30'd231362949;
array2[10503]=30'd231362949;
array2[10504]=30'd231364996;
array2[10505]=30'd228216193;
array2[10506]=30'd228216193;
array2[10507]=30'd231362949;
array2[10508]=30'd231362949;
array2[10509]=30'd231362949;
array2[10510]=30'd231362949;
array2[10511]=30'd231362949;
array2[10512]=30'd231364996;
array2[10513]=30'd231364996;
array2[10514]=30'd231362949;
array2[10515]=30'd234504581;
array2[10516]=30'd231362949;
array2[10517]=30'd231362949;
array2[10518]=30'd231359873;
array2[10519]=30'd231362949;
array2[10520]=30'd231362949;
array2[10521]=30'd229266819;
array2[10522]=30'd231362949;
array2[10523]=30'd231362949;
array2[10524]=30'd231362949;
array2[10525]=30'd231362949;
array2[10526]=30'd231364996;
array2[10527]=30'd229266819;
array2[10528]=30'd231364996;
array2[10529]=30'd231362949;
array2[10530]=30'd231359873;
array2[10531]=30'd231362949;
array2[10532]=30'd231362949;
array2[10533]=30'd231359873;
array2[10534]=30'd231362949;
array2[10535]=30'd231364996;
array2[10536]=30'd229266819;
array2[10537]=30'd234504581;
array2[10538]=30'd231362949;
array2[10539]=30'd234504581;
array2[10540]=30'd231362949;
array2[10541]=30'd231362949;
array2[10542]=30'd229266819;
array2[10543]=30'd231362949;
array2[10544]=30'd231364996;
array2[10545]=30'd231362949;
array2[10546]=30'd272255371;
array2[10547]=30'd532258209;
array2[10548]=30'd272255371;
array2[10549]=30'd230307208;
array2[10550]=30'd234504581;
array2[10551]=30'd231362949;
array2[10552]=30'd230317442;
array2[10553]=30'd229266819;
array2[10554]=30'd228216193;
array2[10555]=30'd228216193;
array2[10556]=30'd231362949;
array2[10557]=30'd231362949;
array2[10558]=30'd230317442;
array2[10559]=30'd231362949;
array2[10560]=30'd212454818;
array2[10561]=30'd234504581;
array2[10562]=30'd228212100;
array2[10563]=30'd231362949;
array2[10564]=30'd229266819;
array2[10565]=30'd229266819;
array2[10566]=30'd229266819;
array2[10567]=30'd231364996;
array2[10568]=30'd229266819;
array2[10569]=30'd229266819;
array2[10570]=30'd231362949;
array2[10571]=30'd229266819;
array2[10572]=30'd231362949;
array2[10573]=30'd234504581;
array2[10574]=30'd231362949;
array2[10575]=30'd231362949;
array2[10576]=30'd231362949;
array2[10577]=30'd231364996;
array2[10578]=30'd230317442;
array2[10579]=30'd231364996;
array2[10580]=30'd231362949;
array2[10581]=30'd231364996;
array2[10582]=30'd231362949;
array2[10583]=30'd231362949;
array2[10584]=30'd229266819;
array2[10585]=30'd228216193;
array2[10586]=30'd231362949;
array2[10587]=30'd231362949;
array2[10588]=30'd231359873;
array2[10589]=30'd231362949;
array2[10590]=30'd231362949;
array2[10591]=30'd231362949;
array2[10592]=30'd231362949;
array2[10593]=30'd229266819;
array2[10594]=30'd231362949;
array2[10595]=30'd229266819;
array2[10596]=30'd230317442;
array2[10597]=30'd229266819;
array2[10598]=30'd231364996;
array2[10599]=30'd229266819;
array2[10600]=30'd231362949;
array2[10601]=30'd229266819;
array2[10602]=30'd229266819;
array2[10603]=30'd231359873;
array2[10604]=30'd231362949;
array2[10605]=30'd231362949;
array2[10606]=30'd231362949;
array2[10607]=30'd229266819;
array2[10608]=30'd230317442;
array2[10609]=30'd231362949;
array2[10610]=30'd231359873;
array2[10611]=30'd228216193;
array2[10612]=30'd229266819;
array2[10613]=30'd230317442;
array2[10614]=30'd229266819;
array2[10615]=30'd228216193;
array2[10616]=30'd230317442;
array2[10617]=30'd230317442;
array2[10618]=30'd230317442;
array2[10619]=30'd231362949;
array2[10620]=30'd231362949;
array2[10621]=30'd231362949;
array2[10622]=30'd231359873;
array2[10623]=30'd229266819;
array2[10624]=30'd228216193;
array2[10625]=30'd230317442;
array2[10626]=30'd230317442;
array2[10627]=30'd230317442;
array2[10628]=30'd231362949;
array2[10629]=30'd229266819;
array2[10630]=30'd231362949;
array2[10631]=30'd228216193;
array2[10632]=30'd231362949;
array2[10633]=30'd231362949;
array2[10634]=30'd229266819;
array2[10635]=30'd231364996;
array2[10636]=30'd231362949;
array2[10637]=30'd231362949;
array2[10638]=30'd231364996;
array2[10639]=30'd231364996;
array2[10640]=30'd231362949;
array2[10641]=30'd229266819;
array2[10642]=30'd234504581;
array2[10643]=30'd230317442;
array2[10644]=30'd229266819;
array2[10645]=30'd231362949;
array2[10646]=30'd231362949;
array2[10647]=30'd234504581;
array2[10648]=30'd231362949;
array2[10649]=30'd231362949;
array2[10650]=30'd230317442;
array2[10651]=30'd231362949;
array2[10652]=30'd229266819;
array2[10653]=30'd231359873;
array2[10654]=30'd231364996;
array2[10655]=30'd230317442;
array2[10656]=30'd212454818;
array2[10657]=30'd234504581;
array2[10658]=30'd228212100;
array2[10659]=30'd230317442;
array2[10660]=30'd231364996;
array2[10661]=30'd231364996;
array2[10662]=30'd231362949;
array2[10663]=30'd231362949;
array2[10664]=30'd228216193;
array2[10665]=30'd229266819;
array2[10666]=30'd229266819;
array2[10667]=30'd231359873;
array2[10668]=30'd231362949;
array2[10669]=30'd231362949;
array2[10670]=30'd231362949;
array2[10671]=30'd231362949;
array2[10672]=30'd230317442;
array2[10673]=30'd231362949;
array2[10674]=30'd229266819;
array2[10675]=30'd228216193;
array2[10676]=30'd229266819;
array2[10677]=30'd230317442;
array2[10678]=30'd231364996;
array2[10679]=30'd231364996;
array2[10680]=30'd231364996;
array2[10681]=30'd231362949;
array2[10682]=30'd231362949;
array2[10683]=30'd229266819;
array2[10684]=30'd228216193;
array2[10685]=30'd229266819;
array2[10686]=30'd231362949;
array2[10687]=30'd231359873;
array2[10688]=30'd231362949;
array2[10689]=30'd231362949;
array2[10690]=30'd231362949;
array2[10691]=30'd231362949;
array2[10692]=30'd229266819;
array2[10693]=30'd231362949;
array2[10694]=30'd229266819;
array2[10695]=30'd229266819;
array2[10696]=30'd230317442;
array2[10697]=30'd230317442;
array2[10698]=30'd231364996;
array2[10699]=30'd231362949;
array2[10700]=30'd230317442;
array2[10701]=30'd231362949;
array2[10702]=30'd231362949;
array2[10703]=30'd228216193;
array2[10704]=30'd231362949;
array2[10705]=30'd231362949;
array2[10706]=30'd231362949;
array2[10707]=30'd231362949;
array2[10708]=30'd231362949;
array2[10709]=30'd231362949;
array2[10710]=30'd231359873;
array2[10711]=30'd230317442;
array2[10712]=30'd230317442;
array2[10713]=30'd231362949;
array2[10714]=30'd229266819;
array2[10715]=30'd231362949;
array2[10716]=30'd230317442;
array2[10717]=30'd231364996;
array2[10718]=30'd230317442;
array2[10719]=30'd230317442;
array2[10720]=30'd231364996;
array2[10721]=30'd231362949;
array2[10722]=30'd231362949;
array2[10723]=30'd231362949;
array2[10724]=30'd228216193;
array2[10725]=30'd229266819;
array2[10726]=30'd229266819;
array2[10727]=30'd231362949;
array2[10728]=30'd229266819;
array2[10729]=30'd231362949;
array2[10730]=30'd231362949;
array2[10731]=30'd230317442;
array2[10732]=30'd230317442;
array2[10733]=30'd231362949;
array2[10734]=30'd229266819;
array2[10735]=30'd231362949;
array2[10736]=30'd230317442;
array2[10737]=30'd231362949;
array2[10738]=30'd231362949;
array2[10739]=30'd230317442;
array2[10740]=30'd229266819;
array2[10741]=30'd229266819;
array2[10742]=30'd229266819;
array2[10743]=30'd228216193;
array2[10744]=30'd231364996;
array2[10745]=30'd230317442;
array2[10746]=30'd229266819;
array2[10747]=30'd229266819;
array2[10748]=30'd231364996;
array2[10749]=30'd231362949;
array2[10750]=30'd231359873;
array2[10751]=30'd231362949;
array2[10752]=30'd193577377;
array2[10753]=30'd227165569;
array2[10754]=30'd228212100;
array2[10755]=30'd231362949;
array2[10756]=30'd231362949;
array2[10757]=30'd231362949;
array2[10758]=30'd231362949;
array2[10759]=30'd231362949;
array2[10760]=30'd231364996;
array2[10761]=30'd231362949;
array2[10762]=30'd229266819;
array2[10763]=30'd231362949;
array2[10764]=30'd231362949;
array2[10765]=30'd234504581;
array2[10766]=30'd231362949;
array2[10767]=30'd231362949;
array2[10768]=30'd229266819;
array2[10769]=30'd231364996;
array2[10770]=30'd231364996;
array2[10771]=30'd231362949;
array2[10772]=30'd231362949;
array2[10773]=30'd231362949;
array2[10774]=30'd231364996;
array2[10775]=30'd231364996;
array2[10776]=30'd231362949;
array2[10777]=30'd230317442;
array2[10778]=30'd231359873;
array2[10779]=30'd229266819;
array2[10780]=30'd231362949;
array2[10781]=30'd231362949;
array2[10782]=30'd231362949;
array2[10783]=30'd231362949;
array2[10784]=30'd234504581;
array2[10785]=30'd229266819;
array2[10786]=30'd231364996;
array2[10787]=30'd231362949;
array2[10788]=30'd231359873;
array2[10789]=30'd228216193;
array2[10790]=30'd234504581;
array2[10791]=30'd230317442;
array2[10792]=30'd231362949;
array2[10793]=30'd227165569;
array2[10794]=30'd229266819;
array2[10795]=30'd231359873;
array2[10796]=30'd231364996;
array2[10797]=30'd230317442;
array2[10798]=30'd229266819;
array2[10799]=30'd229266819;
array2[10800]=30'd234504581;
array2[10801]=30'd231362949;
array2[10802]=30'd231362949;
array2[10803]=30'd231362949;
array2[10804]=30'd231359873;
array2[10805]=30'd229270912;
array2[10806]=30'd231362949;
array2[10807]=30'd231362949;
array2[10808]=30'd231362949;
array2[10809]=30'd234504581;
array2[10810]=30'd231364996;
array2[10811]=30'd231362949;
array2[10812]=30'd230317442;
array2[10813]=30'd230317442;
array2[10814]=30'd231364996;
array2[10815]=30'd231362949;
array2[10816]=30'd231362949;
array2[10817]=30'd228216193;
array2[10818]=30'd229266819;
array2[10819]=30'd229266819;
array2[10820]=30'd231359873;
array2[10821]=30'd231362949;
array2[10822]=30'd234504581;
array2[10823]=30'd231362949;
array2[10824]=30'd231362949;
array2[10825]=30'd230317442;
array2[10826]=30'd231362949;
array2[10827]=30'd229266819;
array2[10828]=30'd228216193;
array2[10829]=30'd230317442;
array2[10830]=30'd230317442;
array2[10831]=30'd229270912;
array2[10832]=30'd230317442;
array2[10833]=30'd228216193;
array2[10834]=30'd234504581;
array2[10835]=30'd228216193;
array2[10836]=30'd234504581;
array2[10837]=30'd234504581;
array2[10838]=30'd229266819;
array2[10839]=30'd231362949;
array2[10840]=30'd231364996;
array2[10841]=30'd229266819;
array2[10842]=30'd228216193;
array2[10843]=30'd229266819;
array2[10844]=30'd231362949;
array2[10845]=30'd229266819;
array2[10846]=30'd231362949;
array2[10847]=30'd231362949;
array2[10848]=30'd338288022;
array2[10849]=30'd272255371;
array2[10850]=30'd227165569;
array2[10851]=30'd231362949;
array2[10852]=30'd229266819;
array2[10853]=30'd231364996;
array2[10854]=30'd225072515;
array2[10855]=30'd228216193;
array2[10856]=30'd231362949;
array2[10857]=30'd228216193;
array2[10858]=30'd229266819;
array2[10859]=30'd229266819;
array2[10860]=30'd231362949;
array2[10861]=30'd231359873;
array2[10862]=30'd231362949;
array2[10863]=30'd231362949;
array2[10864]=30'd231362949;
array2[10865]=30'd230317442;
array2[10866]=30'd229266819;
array2[10867]=30'd231362949;
array2[10868]=30'd228216193;
array2[10869]=30'd229266819;
array2[10870]=30'd230317442;
array2[10871]=30'd229270912;
array2[10872]=30'd256519562;
array2[10873]=30'd227165569;
array2[10874]=30'd234504581;
array2[10875]=30'd229266819;
array2[10876]=30'd229270912;
array2[10877]=30'd229266819;
array2[10878]=30'd229266819;
array2[10879]=30'd231362949;
array2[10880]=30'd230317442;
array2[10881]=30'd231362949;
array2[10882]=30'd231362949;
array2[10883]=30'd231364996;
array2[10884]=30'd231362949;
array2[10885]=30'd231362949;
array2[10886]=30'd231362949;
array2[10887]=30'd228216193;
array2[10888]=30'd230317442;
array2[10889]=30'd229266819;
array2[10890]=30'd231359873;
array2[10891]=30'd231362949;
array2[10892]=30'd231362949;
array2[10893]=30'd231362949;
array2[10894]=30'd231364996;
array2[10895]=30'd230317442;
array2[10896]=30'd234504581;
array2[10897]=30'd229266819;
array2[10898]=30'd231359873;
array2[10899]=30'd230317442;
array2[10900]=30'd230317442;
array2[10901]=30'd230317442;
array2[10902]=30'd230317442;
array2[10903]=30'd228216193;
array2[10904]=30'd234504581;
array2[10905]=30'd231364996;
array2[10906]=30'd231364996;
array2[10907]=30'd231362949;
array2[10908]=30'd229266819;
array2[10909]=30'd229266819;
array2[10910]=30'd228216193;
array2[10911]=30'd229266819;
array2[10912]=30'd229266819;
array2[10913]=30'd231362949;
array2[10914]=30'd231362949;
array2[10915]=30'd231362949;
array2[10916]=30'd231362949;
array2[10917]=30'd231362949;
array2[10918]=30'd230317442;
array2[10919]=30'd231362949;
array2[10920]=30'd229266819;
array2[10921]=30'd228216193;
array2[10922]=30'd230317442;
array2[10923]=30'd230317442;
array2[10924]=30'd230317442;
array2[10925]=30'd230317442;
array2[10926]=30'd231362949;
array2[10927]=30'd234504581;
array2[10928]=30'd231362949;
array2[10929]=30'd231359873;
array2[10930]=30'd231364996;
array2[10931]=30'd229266819;
array2[10932]=30'd228216193;
array2[10933]=30'd231362949;
array2[10934]=30'd231362949;
array2[10935]=30'd231362949;
array2[10936]=30'd231362949;
array2[10937]=30'd229266819;
array2[10938]=30'd231359873;
array2[10939]=30'd231362949;
array2[10940]=30'd231364996;
array2[10941]=30'd231362949;
array2[10942]=30'd229266819;
array2[10943]=30'd231364996;
array2[10944]=30'd304706973;
array2[10945]=30'd377085336;
array2[10946]=30'd377085336;
array2[10947]=30'd229266819;
array2[10948]=30'd231362949;
array2[10949]=30'd401193372;
array2[10950]=30'd603537847;
array2[10951]=30'd272255371;
array2[10952]=30'd227165569;
array2[10953]=30'd229266819;
array2[10954]=30'd229266819;
array2[10955]=30'd230317442;
array2[10956]=30'd230317442;
array2[10957]=30'd229266819;
array2[10958]=30'd231364996;
array2[10959]=30'd229266819;
array2[10960]=30'd228216193;
array2[10961]=30'd220861839;
array2[10962]=30'd221916546;
array2[10963]=30'd234504581;
array2[10964]=30'd231362949;
array2[10965]=30'd234504581;
array2[10966]=30'd231362949;
array2[10967]=30'd231362949;
array2[10968]=30'd338288022;
array2[10969]=30'd377085336;
array2[10970]=30'd236604812;
array2[10971]=30'd231364996;
array2[10972]=30'd256519562;
array2[10973]=30'd603537847;
array2[10974]=30'd377085336;
array2[10975]=30'd231362949;
array2[10976]=30'd231362949;
array2[10977]=30'd231362949;
array2[10978]=30'd230317442;
array2[10979]=30'd229266819;
array2[10980]=30'd231364996;
array2[10981]=30'd231362949;
array2[10982]=30'd229266819;
array2[10983]=30'd229266819;
array2[10984]=30'd229266819;
array2[10985]=30'd231359873;
array2[10986]=30'd231362949;
array2[10987]=30'd231362949;
array2[10988]=30'd231362949;
array2[10989]=30'd231362949;
array2[10990]=30'd231364996;
array2[10991]=30'd229266819;
array2[10992]=30'd231364996;
array2[10993]=30'd229266819;
array2[10994]=30'd231359873;
array2[10995]=30'd229266819;
array2[10996]=30'd231362949;
array2[10997]=30'd229270912;
array2[10998]=30'd230317442;
array2[10999]=30'd229266819;
array2[11000]=30'd228216193;
array2[11001]=30'd229266819;
array2[11002]=30'd234504581;
array2[11003]=30'd231362949;
array2[11004]=30'd231362949;
array2[11005]=30'd231362949;
array2[11006]=30'd229266819;
array2[11007]=30'd231362949;
array2[11008]=30'd229266819;
array2[11009]=30'd229266819;
array2[11010]=30'd229266819;
array2[11011]=30'd231364996;
array2[11012]=30'd230317442;
array2[11013]=30'd231362949;
array2[11014]=30'd231362949;
array2[11015]=30'd228216193;
array2[11016]=30'd230317442;
array2[11017]=30'd229266819;
array2[11018]=30'd228216193;
array2[11019]=30'd231362949;
array2[11020]=30'd231362949;
array2[11021]=30'd231362949;
array2[11022]=30'd231362949;
array2[11023]=30'd231362949;
array2[11024]=30'd231362949;
array2[11025]=30'd231364996;
array2[11026]=30'd228216193;
array2[11027]=30'd231362949;
array2[11028]=30'd229266819;
array2[11029]=30'd231364996;
array2[11030]=30'd230317442;
array2[11031]=30'd229266819;
array2[11032]=30'd234504581;
array2[11033]=30'd229266819;
array2[11034]=30'd234504581;
array2[11035]=30'd230317442;
array2[11036]=30'd230317442;
array2[11037]=30'd231364996;
array2[11038]=30'd231362949;
array2[11039]=30'd231362949;
array2[11040]=30'd338288022;
array2[11041]=30'd338288022;
array2[11042]=30'd272255371;
array2[11043]=30'd228216193;
array2[11044]=30'd228216193;
array2[11045]=30'd377085336;
array2[11046]=30'd532258209;
array2[11047]=30'd272255371;
array2[11048]=30'd227165569;
array2[11049]=30'd229266819;
array2[11050]=30'd227165569;
array2[11051]=30'd231359873;
array2[11052]=30'd231359873;
array2[11053]=30'd231362949;
array2[11054]=30'd230317442;
array2[11055]=30'd229266819;
array2[11056]=30'd227159434;
array2[11057]=30'd208120309;
array2[11058]=30'd179916222;
array2[11059]=30'd228181405;
array2[11060]=30'd213516691;
array2[11061]=30'd213516691;
array2[11062]=30'd234499470;
array2[11063]=30'd231364996;
array2[11064]=30'd301610387;
array2[11065]=30'd301610387;
array2[11066]=30'd236604812;
array2[11067]=30'd231359873;
array2[11068]=30'd256519562;
array2[11069]=30'd553231776;
array2[11070]=30'd338288022;
array2[11071]=30'd231359873;
array2[11072]=30'd234504581;
array2[11073]=30'd231362949;
array2[11074]=30'd229266819;
array2[11075]=30'd231359873;
array2[11076]=30'd234504581;
array2[11077]=30'd231364996;
array2[11078]=30'd231362949;
array2[11079]=30'd229266819;
array2[11080]=30'd231362949;
array2[11081]=30'd229266819;
array2[11082]=30'd231362949;
array2[11083]=30'd231362949;
array2[11084]=30'd234504581;
array2[11085]=30'd231362949;
array2[11086]=30'd231364996;
array2[11087]=30'd231362949;
array2[11088]=30'd231362949;
array2[11089]=30'd231362949;
array2[11090]=30'd231359873;
array2[11091]=30'd231362949;
array2[11092]=30'd231362949;
array2[11093]=30'd230317442;
array2[11094]=30'd228216193;
array2[11095]=30'd231359873;
array2[11096]=30'd231362949;
array2[11097]=30'd231362949;
array2[11098]=30'd228216193;
array2[11099]=30'd231362949;
array2[11100]=30'd231362949;
array2[11101]=30'd231362949;
array2[11102]=30'd231362949;
array2[11103]=30'd228216193;
array2[11104]=30'd229266819;
array2[11105]=30'd231364996;
array2[11106]=30'd231364996;
array2[11107]=30'd231359873;
array2[11108]=30'd229266819;
array2[11109]=30'd231362949;
array2[11110]=30'd231362949;
array2[11111]=30'd229270912;
array2[11112]=30'd229266819;
array2[11113]=30'd228216193;
array2[11114]=30'd231359873;
array2[11115]=30'd231362949;
array2[11116]=30'd231362949;
array2[11117]=30'd229266819;
array2[11118]=30'd229266819;
array2[11119]=30'd231362949;
array2[11120]=30'd229266819;
array2[11121]=30'd230317442;
array2[11122]=30'd231364996;
array2[11123]=30'd231362949;
array2[11124]=30'd229266819;
array2[11125]=30'd231362949;
array2[11126]=30'd231362949;
array2[11127]=30'd229266819;
array2[11128]=30'd229266819;
array2[11129]=30'd231362949;
array2[11130]=30'd231362949;
array2[11131]=30'd228216193;
array2[11132]=30'd229266819;
array2[11133]=30'd229266819;
array2[11134]=30'd229266819;
array2[11135]=30'd231362949;
array2[11136]=30'd304706973;
array2[11137]=30'd256519562;
array2[11138]=30'd227165569;
array2[11139]=30'd228216193;
array2[11140]=30'd231362949;
array2[11141]=30'd228216193;
array2[11142]=30'd228212100;
array2[11143]=30'd227165569;
array2[11144]=30'd234504581;
array2[11145]=30'd234504581;
array2[11146]=30'd229266819;
array2[11147]=30'd229266819;
array2[11148]=30'd231362949;
array2[11149]=30'd228216193;
array2[11150]=30'd228216193;
array2[11151]=30'd231362949;
array2[11152]=30'd281654691;
array2[11153]=30'd407216718;
array2[11154]=30'd444954173;
array2[11155]=30'd444954173;
array2[11156]=30'd444954173;
array2[11157]=30'd407216718;
array2[11158]=30'd260631016;
array2[11159]=30'd228181405;
array2[11160]=30'd248105365;
array2[11161]=30'd230307208;
array2[11162]=30'd231364996;
array2[11163]=30'd231364996;
array2[11164]=30'd229266819;
array2[11165]=30'd225072515;
array2[11166]=30'd230307208;
array2[11167]=30'd234504581;
array2[11168]=30'd229266819;
array2[11169]=30'd231364996;
array2[11170]=30'd231359873;
array2[11171]=30'd231364996;
array2[11172]=30'd231362949;
array2[11173]=30'd229266819;
array2[11174]=30'd231362949;
array2[11175]=30'd231362949;
array2[11176]=30'd231362949;
array2[11177]=30'd229266819;
array2[11178]=30'd231362949;
array2[11179]=30'd230317442;
array2[11180]=30'd231364996;
array2[11181]=30'd231364996;
array2[11182]=30'd231362949;
array2[11183]=30'd234504581;
array2[11184]=30'd231362949;
array2[11185]=30'd231362949;
array2[11186]=30'd229266819;
array2[11187]=30'd229266819;
array2[11188]=30'd228216193;
array2[11189]=30'd231362949;
array2[11190]=30'd231362949;
array2[11191]=30'd231362949;
array2[11192]=30'd231364996;
array2[11193]=30'd229266819;
array2[11194]=30'd229266819;
array2[11195]=30'd231362949;
array2[11196]=30'd231362949;
array2[11197]=30'd231362949;
array2[11198]=30'd231362949;
array2[11199]=30'd231362949;
array2[11200]=30'd231362949;
array2[11201]=30'd229270912;
array2[11202]=30'd231362949;
array2[11203]=30'd231359873;
array2[11204]=30'd228216193;
array2[11205]=30'd231362949;
array2[11206]=30'd230317442;
array2[11207]=30'd231362949;
array2[11208]=30'd229266819;
array2[11209]=30'd231359873;
array2[11210]=30'd231362949;
array2[11211]=30'd231362949;
array2[11212]=30'd230317442;
array2[11213]=30'd231364996;
array2[11214]=30'd229266819;
array2[11215]=30'd228216193;
array2[11216]=30'd231362949;
array2[11217]=30'd229266819;
array2[11218]=30'd230317442;
array2[11219]=30'd231362949;
array2[11220]=30'd231362949;
array2[11221]=30'd234504581;
array2[11222]=30'd231362949;
array2[11223]=30'd231362949;
array2[11224]=30'd229266819;
array2[11225]=30'd231362949;
array2[11226]=30'd229266819;
array2[11227]=30'd229266819;
array2[11228]=30'd230317442;
array2[11229]=30'd230317442;
array2[11230]=30'd230317442;
array2[11231]=30'd231362949;
array2[11232]=30'd212454818;
array2[11233]=30'd234504581;
array2[11234]=30'd227165569;
array2[11235]=30'd229266819;
array2[11236]=30'd230317442;
array2[11237]=30'd230317442;
array2[11238]=30'd230317442;
array2[11239]=30'd231362949;
array2[11240]=30'd231362949;
array2[11241]=30'd229266819;
array2[11242]=30'd231362949;
array2[11243]=30'd230317442;
array2[11244]=30'd229266819;
array2[11245]=30'd231359873;
array2[11246]=30'd231362949;
array2[11247]=30'd234504581;
array2[11248]=30'd281654691;
array2[11249]=30'd560184961;
array2[11250]=30'd799112870;
array2[11251]=30'd828452495;
array2[11252]=30'd828452495;
array2[11253]=30'd768729747;
array2[11254]=30'd538207812;
array2[11255]=30'd483727963;
array2[11256]=30'd319215128;
array2[11257]=30'd193577377;
array2[11258]=30'd212454818;
array2[11259]=30'd227165569;
array2[11260]=30'd231362949;
array2[11261]=30'd231362949;
array2[11262]=30'd230317442;
array2[11263]=30'd229266819;
array2[11264]=30'd229266819;
array2[11265]=30'd231362949;
array2[11266]=30'd234504581;
array2[11267]=30'd231362949;
array2[11268]=30'd231362949;
array2[11269]=30'd231362949;
array2[11270]=30'd231362949;
array2[11271]=30'd231364996;
array2[11272]=30'd231364996;
array2[11273]=30'd229266819;
array2[11274]=30'd231362949;
array2[11275]=30'd231362949;
array2[11276]=30'd230317442;
array2[11277]=30'd231362949;
array2[11278]=30'd229266819;
array2[11279]=30'd231359873;
array2[11280]=30'd231362949;
array2[11281]=30'd231362949;
array2[11282]=30'd230317442;
array2[11283]=30'd230317442;
array2[11284]=30'd231362949;
array2[11285]=30'd231362949;
array2[11286]=30'd231362949;
array2[11287]=30'd228216193;
array2[11288]=30'd229266819;
array2[11289]=30'd229266819;
array2[11290]=30'd231359873;
array2[11291]=30'd231362949;
array2[11292]=30'd231362949;
array2[11293]=30'd231362949;
array2[11294]=30'd231362949;
array2[11295]=30'd229266819;
array2[11296]=30'd231362949;
array2[11297]=30'd229266819;
array2[11298]=30'd229266819;
array2[11299]=30'd230317442;
array2[11300]=30'd230317442;
array2[11301]=30'd231364996;
array2[11302]=30'd229266819;
array2[11303]=30'd228216193;
array2[11304]=30'd234504581;
array2[11305]=30'd231362949;
array2[11306]=30'd231362949;
array2[11307]=30'd231362949;
array2[11308]=30'd231362949;
array2[11309]=30'd231362949;
array2[11310]=30'd231362949;
array2[11311]=30'd229266819;
array2[11312]=30'd230317442;
array2[11313]=30'd231362949;
array2[11314]=30'd229266819;
array2[11315]=30'd229266819;
array2[11316]=30'd229266819;
array2[11317]=30'd231362949;
array2[11318]=30'd231364996;
array2[11319]=30'd229266819;
array2[11320]=30'd228216193;
array2[11321]=30'd231362949;
array2[11322]=30'd231362949;
array2[11323]=30'd230317442;
array2[11324]=30'd229266819;
array2[11325]=30'd231362949;
array2[11326]=30'd231362949;
array2[11327]=30'd231364996;
array2[11328]=30'd193577377;
array2[11329]=30'd227165569;
array2[11330]=30'd228212100;
array2[11331]=30'd231359873;
array2[11332]=30'd230317442;
array2[11333]=30'd230317442;
array2[11334]=30'd231362949;
array2[11335]=30'd231362949;
array2[11336]=30'd231362949;
array2[11337]=30'd228216193;
array2[11338]=30'd229266819;
array2[11339]=30'd231362949;
array2[11340]=30'd231362949;
array2[11341]=30'd229266819;
array2[11342]=30'd231362949;
array2[11343]=30'd234504581;
array2[11344]=30'd232392085;
array2[11345]=30'd538207812;
array2[11346]=30'd851505800;
array2[11347]=30'd851505800;
array2[11348]=30'd851505800;
array2[11349]=30'd858839683;
array2[11350]=30'd851505800;
array2[11351]=30'd828452495;
array2[11352]=30'd727851632;
array2[11353]=30'd645112409;
array2[11354]=30'd560184961;
array2[11355]=30'd179916222;
array2[11356]=30'd179916222;
array2[11357]=30'd193577377;
array2[11358]=30'd231364996;
array2[11359]=30'd231362949;
array2[11360]=30'd231362949;
array2[11361]=30'd231362949;
array2[11362]=30'd231362949;
array2[11363]=30'd231364996;
array2[11364]=30'd229266819;
array2[11365]=30'd231362949;
array2[11366]=30'd231362949;
array2[11367]=30'd231359873;
array2[11368]=30'd231364996;
array2[11369]=30'd229266819;
array2[11370]=30'd229266819;
array2[11371]=30'd231362949;
array2[11372]=30'd231364996;
array2[11373]=30'd234504581;
array2[11374]=30'd231362949;
array2[11375]=30'd231362949;
array2[11376]=30'd234504581;
array2[11377]=30'd229270912;
array2[11378]=30'd231362949;
array2[11379]=30'd228216193;
array2[11380]=30'd231362949;
array2[11381]=30'd231362949;
array2[11382]=30'd231364996;
array2[11383]=30'd231362949;
array2[11384]=30'd228216193;
array2[11385]=30'd229266819;
array2[11386]=30'd229266819;
array2[11387]=30'd231362949;
array2[11388]=30'd231362949;
array2[11389]=30'd231362949;
array2[11390]=30'd231362949;
array2[11391]=30'd231364996;
array2[11392]=30'd231362949;
array2[11393]=30'd228216193;
array2[11394]=30'd231364996;
array2[11395]=30'd231362949;
array2[11396]=30'd231362949;
array2[11397]=30'd231362949;
array2[11398]=30'd234504581;
array2[11399]=30'd230317442;
array2[11400]=30'd231362949;
array2[11401]=30'd229266819;
array2[11402]=30'd231359873;
array2[11403]=30'd231362949;
array2[11404]=30'd231362949;
array2[11405]=30'd231364996;
array2[11406]=30'd231362949;
array2[11407]=30'd231362949;
array2[11408]=30'd228216193;
array2[11409]=30'd231362949;
array2[11410]=30'd231359873;
array2[11411]=30'd229266819;
array2[11412]=30'd231362949;
array2[11413]=30'd231362949;
array2[11414]=30'd231362949;
array2[11415]=30'd231364996;
array2[11416]=30'd229266819;
array2[11417]=30'd229266819;
array2[11418]=30'd231362949;
array2[11419]=30'd231362949;
array2[11420]=30'd229266819;
array2[11421]=30'd229266819;
array2[11422]=30'd228216193;
array2[11423]=30'd231364996;
array2[11424]=30'd212454818;
array2[11425]=30'd234504581;
array2[11426]=30'd228212100;
array2[11427]=30'd230317442;
array2[11428]=30'd230317442;
array2[11429]=30'd230317442;
array2[11430]=30'd231362949;
array2[11431]=30'd230317442;
array2[11432]=30'd229270912;
array2[11433]=30'd231362949;
array2[11434]=30'd231362949;
array2[11435]=30'd228216193;
array2[11436]=30'd228216193;
array2[11437]=30'd229266819;
array2[11438]=30'd231362949;
array2[11439]=30'd231359873;
array2[11440]=30'd221916546;
array2[11441]=30'd483727963;
array2[11442]=30'd865130113;
array2[11443]=30'd851505800;
array2[11444]=30'd851505800;
array2[11445]=30'd858839683;
array2[11446]=30'd858839683;
array2[11447]=30'd858839683;
array2[11448]=30'd858839683;
array2[11449]=30'd858839683;
array2[11450]=30'd828452495;
array2[11451]=30'd708987491;
array2[11452]=30'd678604396;
array2[11453]=30'd506770009;
array2[11454]=30'd179916222;
array2[11455]=30'd212454818;
array2[11456]=30'd227165569;
array2[11457]=30'd228216193;
array2[11458]=30'd231362949;
array2[11459]=30'd231362949;
array2[11460]=30'd231364996;
array2[11461]=30'd229266819;
array2[11462]=30'd229266819;
array2[11463]=30'd228216193;
array2[11464]=30'd231364996;
array2[11465]=30'd231362949;
array2[11466]=30'd229266819;
array2[11467]=30'd231362949;
array2[11468]=30'd229266819;
array2[11469]=30'd231362949;
array2[11470]=30'd231362949;
array2[11471]=30'd231362949;
array2[11472]=30'd231362949;
array2[11473]=30'd231362949;
array2[11474]=30'd231364996;
array2[11475]=30'd229266819;
array2[11476]=30'd229266819;
array2[11477]=30'd229266819;
array2[11478]=30'd231362949;
array2[11479]=30'd234504581;
array2[11480]=30'd230317442;
array2[11481]=30'd231362949;
array2[11482]=30'd231362949;
array2[11483]=30'd229266819;
array2[11484]=30'd228216193;
array2[11485]=30'd229266819;
array2[11486]=30'd229266819;
array2[11487]=30'd231364996;
array2[11488]=30'd230317442;
array2[11489]=30'd229266819;
array2[11490]=30'd231362949;
array2[11491]=30'd231359873;
array2[11492]=30'd234504581;
array2[11493]=30'd231362949;
array2[11494]=30'd229266819;
array2[11495]=30'd229266819;
array2[11496]=30'd229266819;
array2[11497]=30'd229270912;
array2[11498]=30'd229266819;
array2[11499]=30'd230317442;
array2[11500]=30'd229266819;
array2[11501]=30'd229266819;
array2[11502]=30'd231362949;
array2[11503]=30'd231362949;
array2[11504]=30'd231364996;
array2[11505]=30'd231362949;
array2[11506]=30'd231362949;
array2[11507]=30'd231362949;
array2[11508]=30'd229266819;
array2[11509]=30'd229266819;
array2[11510]=30'd231362949;
array2[11511]=30'd231362949;
array2[11512]=30'd231362949;
array2[11513]=30'd231362949;
array2[11514]=30'd231362949;
array2[11515]=30'd229266819;
array2[11516]=30'd231362949;
array2[11517]=30'd229266819;
array2[11518]=30'd228216193;
array2[11519]=30'd229266819;
array2[11520]=30'd212454818;
array2[11521]=30'd234504581;
array2[11522]=30'd227165569;
array2[11523]=30'd231359873;
array2[11524]=30'd230317442;
array2[11525]=30'd230317442;
array2[11526]=30'd231362949;
array2[11527]=30'd229266819;
array2[11528]=30'd234504581;
array2[11529]=30'd231362949;
array2[11530]=30'd229266819;
array2[11531]=30'd229266819;
array2[11532]=30'd231362949;
array2[11533]=30'd229266819;
array2[11534]=30'd231362949;
array2[11535]=30'd231362949;
array2[11536]=30'd221916546;
array2[11537]=30'd483727963;
array2[11538]=30'd865130113;
array2[11539]=30'd858839683;
array2[11540]=30'd851505800;
array2[11541]=30'd858839683;
array2[11542]=30'd858839683;
array2[11543]=30'd858839683;
array2[11544]=30'd851505800;
array2[11545]=30'd858839683;
array2[11546]=30'd858839683;
array2[11547]=30'd851505800;
array2[11548]=30'd858839683;
array2[11549]=30'd768729747;
array2[11550]=30'd518272648;
array2[11551]=30'd193577377;
array2[11552]=30'd229270912;
array2[11553]=30'd230317442;
array2[11554]=30'd231362949;
array2[11555]=30'd231362949;
array2[11556]=30'd231364996;
array2[11557]=30'd228216193;
array2[11558]=30'd229266819;
array2[11559]=30'd231362949;
array2[11560]=30'd231359873;
array2[11561]=30'd231362949;
array2[11562]=30'd231362949;
array2[11563]=30'd231362949;
array2[11564]=30'd231362949;
array2[11565]=30'd231364996;
array2[11566]=30'd231364996;
array2[11567]=30'd231362949;
array2[11568]=30'd228216193;
array2[11569]=30'd231362949;
array2[11570]=30'd230317442;
array2[11571]=30'd231364996;
array2[11572]=30'd229266819;
array2[11573]=30'd228216193;
array2[11574]=30'd234504581;
array2[11575]=30'd231362949;
array2[11576]=30'd231362949;
array2[11577]=30'd231362949;
array2[11578]=30'd231362949;
array2[11579]=30'd229266819;
array2[11580]=30'd231362949;
array2[11581]=30'd231362949;
array2[11582]=30'd229266819;
array2[11583]=30'd230317442;
array2[11584]=30'd229266819;
array2[11585]=30'd229266819;
array2[11586]=30'd229266819;
array2[11587]=30'd229266819;
array2[11588]=30'd231362949;
array2[11589]=30'd231362949;
array2[11590]=30'd231362949;
array2[11591]=30'd231362949;
array2[11592]=30'd231362949;
array2[11593]=30'd230317442;
array2[11594]=30'd230317442;
array2[11595]=30'd230317442;
array2[11596]=30'd229266819;
array2[11597]=30'd231362949;
array2[11598]=30'd228216193;
array2[11599]=30'd230317442;
array2[11600]=30'd230317442;
array2[11601]=30'd231364996;
array2[11602]=30'd231362949;
array2[11603]=30'd231362949;
array2[11604]=30'd228216193;
array2[11605]=30'd231362949;
array2[11606]=30'd229266819;
array2[11607]=30'd231362949;
array2[11608]=30'd231362949;
array2[11609]=30'd231359873;
array2[11610]=30'd231362949;
array2[11611]=30'd231362949;
array2[11612]=30'd230317442;
array2[11613]=30'd231364996;
array2[11614]=30'd230317442;
array2[11615]=30'd227165569;
array2[11616]=30'd212454818;
array2[11617]=30'd234504581;
array2[11618]=30'd228212100;
array2[11619]=30'd230317442;
array2[11620]=30'd230317442;
array2[11621]=30'd230317442;
array2[11622]=30'd231362949;
array2[11623]=30'd230317442;
array2[11624]=30'd231364996;
array2[11625]=30'd231362949;
array2[11626]=30'd231362949;
array2[11627]=30'd231362949;
array2[11628]=30'd229266819;
array2[11629]=30'd228216193;
array2[11630]=30'd229266819;
array2[11631]=30'd229266819;
array2[11632]=30'd221916546;
array2[11633]=30'd483727963;
array2[11634]=30'd865130113;
array2[11635]=30'd851505800;
array2[11636]=30'd858839683;
array2[11637]=30'd851505800;
array2[11638]=30'd851505800;
array2[11639]=30'd858839683;
array2[11640]=30'd858839683;
array2[11641]=30'd851505800;
array2[11642]=30'd851505800;
array2[11643]=30'd858839683;
array2[11644]=30'd851505800;
array2[11645]=30'd851505800;
array2[11646]=30'd645112409;
array2[11647]=30'd186252693;
array2[11648]=30'd229266819;
array2[11649]=30'd231364996;
array2[11650]=30'd229266819;
array2[11651]=30'd231362949;
array2[11652]=30'd229266819;
array2[11653]=30'd230317442;
array2[11654]=30'd229266819;
array2[11655]=30'd231362949;
array2[11656]=30'd231362949;
array2[11657]=30'd231362949;
array2[11658]=30'd231362949;
array2[11659]=30'd231359873;
array2[11660]=30'd231362949;
array2[11661]=30'd231364996;
array2[11662]=30'd231364996;
array2[11663]=30'd231362949;
array2[11664]=30'd229266819;
array2[11665]=30'd231362949;
array2[11666]=30'd231364996;
array2[11667]=30'd231362949;
array2[11668]=30'd229266819;
array2[11669]=30'd228216193;
array2[11670]=30'd234504581;
array2[11671]=30'd231362949;
array2[11672]=30'd230317442;
array2[11673]=30'd231362949;
array2[11674]=30'd234504581;
array2[11675]=30'd228216193;
array2[11676]=30'd228216193;
array2[11677]=30'd229266819;
array2[11678]=30'd231364996;
array2[11679]=30'd231362949;
array2[11680]=30'd227165569;
array2[11681]=30'd228216193;
array2[11682]=30'd231362949;
array2[11683]=30'd234504581;
array2[11684]=30'd231364996;
array2[11685]=30'd230317442;
array2[11686]=30'd229266819;
array2[11687]=30'd231362949;
array2[11688]=30'd231362949;
array2[11689]=30'd228216193;
array2[11690]=30'd229266819;
array2[11691]=30'd231362949;
array2[11692]=30'd231359873;
array2[11693]=30'd231364996;
array2[11694]=30'd231362949;
array2[11695]=30'd234504581;
array2[11696]=30'd231362949;
array2[11697]=30'd231362949;
array2[11698]=30'd231364996;
array2[11699]=30'd229266819;
array2[11700]=30'd229266819;
array2[11701]=30'd229266819;
array2[11702]=30'd231364996;
array2[11703]=30'd231364996;
array2[11704]=30'd230317442;
array2[11705]=30'd234504581;
array2[11706]=30'd231362949;
array2[11707]=30'd231362949;
array2[11708]=30'd231362949;
array2[11709]=30'd231364996;
array2[11710]=30'd230317442;
array2[11711]=30'd229266819;
array2[11712]=30'd212454818;
array2[11713]=30'd234504581;
array2[11714]=30'd228212100;
array2[11715]=30'd230317442;
array2[11716]=30'd230317442;
array2[11717]=30'd230317442;
array2[11718]=30'd231362949;
array2[11719]=30'd230317442;
array2[11720]=30'd231362949;
array2[11721]=30'd231362949;
array2[11722]=30'd234504581;
array2[11723]=30'd231364996;
array2[11724]=30'd229266819;
array2[11725]=30'd228216193;
array2[11726]=30'd231362949;
array2[11727]=30'd231362949;
array2[11728]=30'd221916546;
array2[11729]=30'd444954173;
array2[11730]=30'd770812573;
array2[11731]=30'd851505800;
array2[11732]=30'd858839683;
array2[11733]=30'd858839683;
array2[11734]=30'd858839683;
array2[11735]=30'd858839683;
array2[11736]=30'd858839683;
array2[11737]=30'd858839683;
array2[11738]=30'd851505800;
array2[11739]=30'd858839683;
array2[11740]=30'd858839683;
array2[11741]=30'd858839683;
array2[11742]=30'd645112409;
array2[11743]=30'd186252693;
array2[11744]=30'd234504581;
array2[11745]=30'd228216193;
array2[11746]=30'd231362949;
array2[11747]=30'd231362949;
array2[11748]=30'd231362949;
array2[11749]=30'd228216193;
array2[11750]=30'd229266819;
array2[11751]=30'd230317442;
array2[11752]=30'd228216193;
array2[11753]=30'd228216193;
array2[11754]=30'd229266819;
array2[11755]=30'd231362949;
array2[11756]=30'd231362949;
array2[11757]=30'd234504581;
array2[11758]=30'd231362949;
array2[11759]=30'd234504581;
array2[11760]=30'd231362949;
array2[11761]=30'd231362949;
array2[11762]=30'd228216193;
array2[11763]=30'd231359873;
array2[11764]=30'd231364996;
array2[11765]=30'd231362949;
array2[11766]=30'd220861839;
array2[11767]=30'd212454818;
array2[11768]=30'd212454818;
array2[11769]=30'd212454818;
array2[11770]=30'd234499470;
array2[11771]=30'd238691720;
array2[11772]=30'd234504581;
array2[11773]=30'd227165569;
array2[11774]=30'd238691720;
array2[11775]=30'd238691720;
array2[11776]=30'd262793620;
array2[11777]=30'd234504581;
array2[11778]=30'd231362949;
array2[11779]=30'd231362949;
array2[11780]=30'd234504581;
array2[11781]=30'd234504581;
array2[11782]=30'd231364996;
array2[11783]=30'd229266819;
array2[11784]=30'd229266819;
array2[11785]=30'd231362949;
array2[11786]=30'd231362949;
array2[11787]=30'd231362949;
array2[11788]=30'd231362949;
array2[11789]=30'd231362949;
array2[11790]=30'd231362949;
array2[11791]=30'd229270912;
array2[11792]=30'd231364996;
array2[11793]=30'd234504581;
array2[11794]=30'd231362949;
array2[11795]=30'd234504581;
array2[11796]=30'd231364996;
array2[11797]=30'd230317442;
array2[11798]=30'd228216193;
array2[11799]=30'd228216193;
array2[11800]=30'd231362949;
array2[11801]=30'd231362949;
array2[11802]=30'd231364996;
array2[11803]=30'd231362949;
array2[11804]=30'd234504581;
array2[11805]=30'd228216193;
array2[11806]=30'd227165569;
array2[11807]=30'd227165569;
array2[11808]=30'd212454818;
array2[11809]=30'd234504581;
array2[11810]=30'd228212100;
array2[11811]=30'd230317442;
array2[11812]=30'd230317442;
array2[11813]=30'd230317442;
array2[11814]=30'd231362949;
array2[11815]=30'd230317442;
array2[11816]=30'd231362949;
array2[11817]=30'd231362949;
array2[11818]=30'd231362949;
array2[11819]=30'd231359873;
array2[11820]=30'd229266819;
array2[11821]=30'd228216193;
array2[11822]=30'd230317442;
array2[11823]=30'd256519562;
array2[11824]=30'd256519562;
array2[11825]=30'd347490866;
array2[11826]=30'd565444213;
array2[11827]=30'd645112409;
array2[11828]=30'd645112409;
array2[11829]=30'd645112409;
array2[11830]=30'd645112409;
array2[11831]=30'd708987491;
array2[11832]=30'd819020415;
array2[11833]=30'd828452495;
array2[11834]=30'd828452495;
array2[11835]=30'd828452495;
array2[11836]=30'd858839683;
array2[11837]=30'd851505800;
array2[11838]=30'd645112409;
array2[11839]=30'd186252693;
array2[11840]=30'd227165569;
array2[11841]=30'd228216193;
array2[11842]=30'd229266819;
array2[11843]=30'd231362949;
array2[11844]=30'd229266819;
array2[11845]=30'd228216193;
array2[11846]=30'd256519562;
array2[11847]=30'd272255371;
array2[11848]=30'd228216193;
array2[11849]=30'd234504581;
array2[11850]=30'd229266819;
array2[11851]=30'd229266819;
array2[11852]=30'd231359873;
array2[11853]=30'd234504581;
array2[11854]=30'd229266819;
array2[11855]=30'd231362949;
array2[11856]=30'd228216193;
array2[11857]=30'd231362949;
array2[11858]=30'd256519562;
array2[11859]=30'd377085336;
array2[11860]=30'd256519562;
array2[11861]=30'd231362949;
array2[11862]=30'd212454818;
array2[11863]=30'd150539724;
array2[11864]=30'd124307934;
array2[11865]=30'd124307934;
array2[11866]=30'd195647926;
array2[11867]=30'd254365107;
array2[11868]=30'd207191473;
array2[11869]=30'd248105365;
array2[11870]=30'd262793620;
array2[11871]=30'd238691720;
array2[11872]=30'd238691720;
array2[11873]=30'd262793620;
array2[11874]=30'd262793620;
array2[11875]=30'd238691720;
array2[11876]=30'd238691720;
array2[11877]=30'd238691720;
array2[11878]=30'd227165569;
array2[11879]=30'd234504581;
array2[11880]=30'd229266819;
array2[11881]=30'd229270912;
array2[11882]=30'd231362949;
array2[11883]=30'd227165569;
array2[11884]=30'd231359873;
array2[11885]=30'd231364996;
array2[11886]=30'd229266819;
array2[11887]=30'd229266819;
array2[11888]=30'd231359873;
array2[11889]=30'd231362949;
array2[11890]=30'd231362949;
array2[11891]=30'd231362949;
array2[11892]=30'd231362949;
array2[11893]=30'd229266819;
array2[11894]=30'd231364996;
array2[11895]=30'd229266819;
array2[11896]=30'd231359873;
array2[11897]=30'd229266819;
array2[11898]=30'd231362949;
array2[11899]=30'd230317442;
array2[11900]=30'd230317442;
array2[11901]=30'd227165569;
array2[11902]=30'd229266819;
array2[11903]=30'd231362949;
array2[11904]=30'd193577377;
array2[11905]=30'd227165569;
array2[11906]=30'd228212100;
array2[11907]=30'd231362949;
array2[11908]=30'd231362949;
array2[11909]=30'd230317442;
array2[11910]=30'd229266819;
array2[11911]=30'd229266819;
array2[11912]=30'd231362949;
array2[11913]=30'd231362949;
array2[11914]=30'd231362949;
array2[11915]=30'd229266819;
array2[11916]=30'd231362949;
array2[11917]=30'd231362949;
array2[11918]=30'd231364996;
array2[11919]=30'd377085336;
array2[11920]=30'd405404052;
array2[11921]=30'd213516691;
array2[11922]=30'd193577377;
array2[11923]=30'd193577377;
array2[11924]=30'd193577377;
array2[11925]=30'd193577377;
array2[11926]=30'd193577377;
array2[11927]=30'd284737060;
array2[11928]=30'd506770009;
array2[11929]=30'd538207812;
array2[11930]=30'd538207812;
array2[11931]=30'd566515308;
array2[11932]=30'd819020415;
array2[11933]=30'd828452495;
array2[11934]=30'd566515308;
array2[11935]=30'd193577377;
array2[11936]=30'd234504581;
array2[11937]=30'd231362949;
array2[11938]=30'd230317442;
array2[11939]=30'd229266819;
array2[11940]=30'd229266819;
array2[11941]=30'd231359873;
array2[11942]=30'd338288022;
array2[11943]=30'd405404052;
array2[11944]=30'd238691720;
array2[11945]=30'd231359873;
array2[11946]=30'd231359873;
array2[11947]=30'd230317442;
array2[11948]=30'd229266819;
array2[11949]=30'd229266819;
array2[11950]=30'd231362949;
array2[11951]=30'd231364996;
array2[11952]=30'd338288022;
array2[11953]=30'd272255371;
array2[11954]=30'd377085336;
array2[11955]=30'd719920570;
array2[11956]=30'd401193372;
array2[11957]=30'd256519562;
array2[11958]=30'd338288022;
array2[11959]=30'd212454818;
array2[11960]=30'd150539724;
array2[11961]=30'd106464746;
array2[11962]=30'd131612152;
array2[11963]=30'd299264555;
array2[11964]=30'd357913199;
array2[11965]=30'd281508345;
array2[11966]=30'd260631016;
array2[11967]=30'd207191473;
array2[11968]=30'd240774546;
array2[11969]=30'd262793620;
array2[11970]=30'd262793620;
array2[11971]=30'd262793620;
array2[11972]=30'd262793620;
array2[11973]=30'd238691720;
array2[11974]=30'd238691720;
array2[11975]=30'd238691720;
array2[11976]=30'd234504581;
array2[11977]=30'd231364996;
array2[11978]=30'd231364996;
array2[11979]=30'd228216193;
array2[11980]=30'd228216193;
array2[11981]=30'd229266819;
array2[11982]=30'd229266819;
array2[11983]=30'd228216193;
array2[11984]=30'd231362949;
array2[11985]=30'd231362949;
array2[11986]=30'd231362949;
array2[11987]=30'd231362949;
array2[11988]=30'd229266819;
array2[11989]=30'd231362949;
array2[11990]=30'd231362949;
array2[11991]=30'd229266819;
array2[11992]=30'd229266819;
array2[11993]=30'd230317442;
array2[11994]=30'd230317442;
array2[11995]=30'd230317442;
array2[11996]=30'd229266819;
array2[11997]=30'd234504581;
array2[11998]=30'd231362949;
array2[11999]=30'd231362949;
array2[12000]=30'd212454818;
array2[12001]=30'd234504581;
array2[12002]=30'd228212100;
array2[12003]=30'd230317442;
array2[12004]=30'd230317442;
array2[12005]=30'd230317442;
array2[12006]=30'd231362949;
array2[12007]=30'd230317442;
array2[12008]=30'd231362949;
array2[12009]=30'd231362949;
array2[12010]=30'd231362949;
array2[12011]=30'd231362949;
array2[12012]=30'd234504581;
array2[12013]=30'd231362949;
array2[12014]=30'd229266819;
array2[12015]=30'd229266819;
array2[12016]=30'd231362949;
array2[12017]=30'd231362949;
array2[12018]=30'd231362949;
array2[12019]=30'd231362949;
array2[12020]=30'd231362949;
array2[12021]=30'd231362949;
array2[12022]=30'd231364996;
array2[12023]=30'd228212100;
array2[12024]=30'd213516691;
array2[12025]=30'd213516691;
array2[12026]=30'd212454818;
array2[12027]=30'd208120309;
array2[12028]=30'd819020415;
array2[12029]=30'd764529268;
array2[12030]=30'd401997362;
array2[12031]=30'd186252693;
array2[12032]=30'd228216193;
array2[12033]=30'd227165569;
array2[12034]=30'd228216193;
array2[12035]=30'd231362949;
array2[12036]=30'd231362949;
array2[12037]=30'd231362949;
array2[12038]=30'd231364996;
array2[12039]=30'd231362949;
array2[12040]=30'd231362949;
array2[12041]=30'd231362949;
array2[12042]=30'd229266819;
array2[12043]=30'd229266819;
array2[12044]=30'd231364996;
array2[12045]=30'd231359873;
array2[12046]=30'd234504581;
array2[12047]=30'd256519562;
array2[12048]=30'd603537847;
array2[12049]=30'd425297329;
array2[12050]=30'd230307208;
array2[12051]=30'd238691720;
array2[12052]=30'd234499470;
array2[12053]=30'd401193372;
array2[12054]=30'd603537847;
array2[12055]=30'd220861839;
array2[12056]=30'd212454818;
array2[12057]=30'd124307934;
array2[12058]=30'd159912438;
array2[12059]=30'd357913199;
array2[12060]=30'd539218630;
array2[12061]=30'd560184961;
array2[12062]=30'd518272648;
array2[12063]=30'd434416250;
array2[12064]=30'd190356956;
array2[12065]=30'd260631016;
array2[12066]=30'd265928088;
array2[12067]=30'd262793620;
array2[12068]=30'd262793620;
array2[12069]=30'd262793620;
array2[12070]=30'd234504581;
array2[12071]=30'd238691720;
array2[12072]=30'd238691720;
array2[12073]=30'd262793620;
array2[12074]=30'd238691720;
array2[12075]=30'd238691720;
array2[12076]=30'd234504581;
array2[12077]=30'd234504581;
array2[12078]=30'd231359873;
array2[12079]=30'd230317442;
array2[12080]=30'd231362949;
array2[12081]=30'd227165569;
array2[12082]=30'd231362949;
array2[12083]=30'd231362949;
array2[12084]=30'd229266819;
array2[12085]=30'd229266819;
array2[12086]=30'd231364996;
array2[12087]=30'd229266819;
array2[12088]=30'd231359873;
array2[12089]=30'd231362949;
array2[12090]=30'd230317442;
array2[12091]=30'd229266819;
array2[12092]=30'd231362949;
array2[12093]=30'd231362949;
array2[12094]=30'd231362949;
array2[12095]=30'd231362949;
array2[12096]=30'd212454818;
array2[12097]=30'd234504581;
array2[12098]=30'd228212100;
array2[12099]=30'd230317442;
array2[12100]=30'd230317442;
array2[12101]=30'd230317442;
array2[12102]=30'd231362949;
array2[12103]=30'd230317442;
array2[12104]=30'd231362949;
array2[12105]=30'd231362949;
array2[12106]=30'd231362949;
array2[12107]=30'd256519562;
array2[12108]=30'd256519562;
array2[12109]=30'd231364996;
array2[12110]=30'd229266819;
array2[12111]=30'd229266819;
array2[12112]=30'd228216193;
array2[12113]=30'd230317442;
array2[12114]=30'd230317442;
array2[12115]=30'd256519562;
array2[12116]=30'd256519562;
array2[12117]=30'd231364996;
array2[12118]=30'd231362949;
array2[12119]=30'd256519562;
array2[12120]=30'd256519562;
array2[12121]=30'd227165569;
array2[12122]=30'd231364996;
array2[12123]=30'd249001484;
array2[12124]=30'd819020415;
array2[12125]=30'd678604396;
array2[12126]=30'd179916222;
array2[12127]=30'd240774546;
array2[12128]=30'd238691720;
array2[12129]=30'd238691720;
array2[12130]=30'd256519562;
array2[12131]=30'd256519562;
array2[12132]=30'd234504581;
array2[12133]=30'd231362949;
array2[12134]=30'd230317442;
array2[12135]=30'd230317442;
array2[12136]=30'd231362949;
array2[12137]=30'd231362949;
array2[12138]=30'd256519562;
array2[12139]=30'd272255371;
array2[12140]=30'd231364996;
array2[12141]=30'd231362949;
array2[12142]=30'd256519562;
array2[12143]=30'd338288022;
array2[12144]=30'd256519562;
array2[12145]=30'd227165569;
array2[12146]=30'd227165569;
array2[12147]=30'd195647926;
array2[12148]=30'd150539724;
array2[12149]=30'd150539724;
array2[12150]=30'd150539724;
array2[12151]=30'd150539724;
array2[12152]=30'd190356956;
array2[12153]=30'd444954173;
array2[12154]=30'd450208341;
array2[12155]=30'd483727963;
array2[12156]=30'd518272648;
array2[12157]=30'd606320275;
array2[12158]=30'd604201637;
array2[12159]=30'd560184961;
array2[12160]=30'd518272648;
array2[12161]=30'd375721588;
array2[12162]=30'd281508345;
array2[12163]=30'd260631016;
array2[12164]=30'd262793620;
array2[12165]=30'd262793620;
array2[12166]=30'd262793620;
array2[12167]=30'd262793620;
array2[12168]=30'd238691720;
array2[12169]=30'd262793620;
array2[12170]=30'd262793620;
array2[12171]=30'd238691720;
array2[12172]=30'd262793620;
array2[12173]=30'd238691720;
array2[12174]=30'd234504581;
array2[12175]=30'd231364996;
array2[12176]=30'd229266819;
array2[12177]=30'd231362949;
array2[12178]=30'd229266819;
array2[12179]=30'd229270912;
array2[12180]=30'd231362949;
array2[12181]=30'd231362949;
array2[12182]=30'd231362949;
array2[12183]=30'd228216193;
array2[12184]=30'd229266819;
array2[12185]=30'd231362949;
array2[12186]=30'd231359873;
array2[12187]=30'd231362949;
array2[12188]=30'd231362949;
array2[12189]=30'd231362949;
array2[12190]=30'd229266819;
array2[12191]=30'd230317442;
array2[12192]=30'd193577377;
array2[12193]=30'd227165569;
array2[12194]=30'd228212100;
array2[12195]=30'd231362949;
array2[12196]=30'd231362949;
array2[12197]=30'd231362949;
array2[12198]=30'd231362949;
array2[12199]=30'd230317442;
array2[12200]=30'd231364996;
array2[12201]=30'd228216193;
array2[12202]=30'd228216193;
array2[12203]=30'd405404052;
array2[12204]=30'd377085336;
array2[12205]=30'd234504581;
array2[12206]=30'd231362949;
array2[12207]=30'd230317442;
array2[12208]=30'd230317442;
array2[12209]=30'd229266819;
array2[12210]=30'd231362949;
array2[12211]=30'd377085336;
array2[12212]=30'd405404052;
array2[12213]=30'd256519562;
array2[12214]=30'd234499470;
array2[12215]=30'd532258209;
array2[12216]=30'd425297329;
array2[12217]=30'd227159434;
array2[12218]=30'd228216193;
array2[12219]=30'd249001484;
array2[12220]=30'd823228019;
array2[12221]=30'd708987491;
array2[12222]=30'd281508345;
array2[12223]=30'd228181405;
array2[12224]=30'd228181405;
array2[12225]=30'd228181405;
array2[12226]=30'd338288022;
array2[12227]=30'd401193372;
array2[12228]=30'd238691720;
array2[12229]=30'd228216193;
array2[12230]=30'd230317442;
array2[12231]=30'd230317442;
array2[12232]=30'd229266819;
array2[12233]=30'd231362949;
array2[12234]=30'd301610387;
array2[12235]=30'd405404052;
array2[12236]=30'd236604812;
array2[12237]=30'd234504581;
array2[12238]=30'd425297329;
array2[12239]=30'd664345022;
array2[12240]=30'd338288022;
array2[12241]=30'd228212100;
array2[12242]=30'd234504581;
array2[12243]=30'd220861839;
array2[12244]=30'd150539724;
array2[12245]=30'd124307934;
array2[12246]=30'd124307934;
array2[12247]=30'd124307934;
array2[12248]=30'd218607140;
array2[12249]=30'd678602388;
array2[12250]=30'd768729747;
array2[12251]=30'd805398138;
array2[12252]=30'd764529268;
array2[12253]=30'd565444213;
array2[12254]=30'd566515308;
array2[12255]=30'd566515308;
array2[12256]=30'd560184961;
array2[12257]=30'd539218630;
array2[12258]=30'd518272648;
array2[12259]=30'd347490866;
array2[12260]=30'd254365107;
array2[12261]=30'd228181405;
array2[12262]=30'd257539480;
array2[12263]=30'd228181405;
array2[12264]=30'd248105365;
array2[12265]=30'd262793620;
array2[12266]=30'd262793620;
array2[12267]=30'd262793620;
array2[12268]=30'd262793620;
array2[12269]=30'd262793620;
array2[12270]=30'd262793620;
array2[12271]=30'd238691720;
array2[12272]=30'd228216193;
array2[12273]=30'd231362949;
array2[12274]=30'd231364996;
array2[12275]=30'd231364996;
array2[12276]=30'd231362949;
array2[12277]=30'd231362949;
array2[12278]=30'd228216193;
array2[12279]=30'd229266819;
array2[12280]=30'd231362949;
array2[12281]=30'd231359873;
array2[12282]=30'd231362949;
array2[12283]=30'd231362949;
array2[12284]=30'd231362949;
array2[12285]=30'd231362949;
array2[12286]=30'd229266819;
array2[12287]=30'd231362949;
array2[12288]=30'd193577377;
array2[12289]=30'd227165569;
array2[12290]=30'd228212100;
array2[12291]=30'd231362949;
array2[12292]=30'd231362949;
array2[12293]=30'd231362949;
array2[12294]=30'd231364996;
array2[12295]=30'd229266819;
array2[12296]=30'd229266819;
array2[12297]=30'd231362949;
array2[12298]=30'd231362949;
array2[12299]=30'd256519562;
array2[12300]=30'd256519562;
array2[12301]=30'd228216193;
array2[12302]=30'd229266819;
array2[12303]=30'd231364996;
array2[12304]=30'd231364996;
array2[12305]=30'd231359873;
array2[12306]=30'd228216193;
array2[12307]=30'd256519562;
array2[12308]=30'd256519562;
array2[12309]=30'd231362949;
array2[12310]=30'd228216193;
array2[12311]=30'd256519562;
array2[12312]=30'd256519562;
array2[12313]=30'd231362949;
array2[12314]=30'd231362949;
array2[12315]=30'd249001484;
array2[12316]=30'd823228019;
array2[12317]=30'd819020415;
array2[12318]=30'd646130287;
array2[12319]=30'd444954173;
array2[12320]=30'd444954173;
array2[12321]=30'd401997362;
array2[12322]=30'd190356956;
array2[12323]=30'd262793620;
array2[12324]=30'd234504581;
array2[12325]=30'd230317442;
array2[12326]=30'd229266819;
array2[12327]=30'd231364996;
array2[12328]=30'd231364996;
array2[12329]=30'd231362949;
array2[12330]=30'd229270912;
array2[12331]=30'd256519562;
array2[12332]=30'd234504581;
array2[12333]=30'd231362949;
array2[12334]=30'd256519562;
array2[12335]=30'd272255371;
array2[12336]=30'd256519562;
array2[12337]=30'd227165569;
array2[12338]=30'd230317442;
array2[12339]=30'd230317442;
array2[12340]=30'd220861839;
array2[12341]=30'd179916222;
array2[12342]=30'd150539724;
array2[12343]=30'd124307934;
array2[12344]=30'd218607140;
array2[12345]=30'd631447172;
array2[12346]=30'd768729747;
array2[12347]=30'd819020415;
array2[12348]=30'd819020415;
array2[12349]=30'd805398138;
array2[12350]=30'd819020415;
array2[12351]=30'd770816666;
array2[12352]=30'd711090860;
array2[12353]=30'd565444213;
array2[12354]=30'd506770009;
array2[12355]=30'd506770009;
array2[12356]=30'd407216718;
array2[12357]=30'd444954173;
array2[12358]=30'd444954173;
array2[12359]=30'd444954173;
array2[12360]=30'd444954173;
array2[12361]=30'd260631016;
array2[12362]=30'd228181405;
array2[12363]=30'd281654691;
array2[12364]=30'd262793620;
array2[12365]=30'd265928088;
array2[12366]=30'd262793620;
array2[12367]=30'd262793620;
array2[12368]=30'd238691720;
array2[12369]=30'd234504581;
array2[12370]=30'd234504581;
array2[12371]=30'd231362949;
array2[12372]=30'd229266819;
array2[12373]=30'd229266819;
array2[12374]=30'd231362949;
array2[12375]=30'd231362949;
array2[12376]=30'd231362949;
array2[12377]=30'd231362949;
array2[12378]=30'd231362949;
array2[12379]=30'd231362949;
array2[12380]=30'd231364996;
array2[12381]=30'd231364996;
array2[12382]=30'd234504581;
array2[12383]=30'd229266819;
array2[12384]=30'd193577377;
array2[12385]=30'd227165569;
array2[12386]=30'd228212100;
array2[12387]=30'd231362949;
array2[12388]=30'd231362949;
array2[12389]=30'd231362949;
array2[12390]=30'd231362949;
array2[12391]=30'd229266819;
array2[12392]=30'd231364996;
array2[12393]=30'd231362949;
array2[12394]=30'd228216193;
array2[12395]=30'd231362949;
array2[12396]=30'd231362949;
array2[12397]=30'd229266819;
array2[12398]=30'd231364996;
array2[12399]=30'd256519562;
array2[12400]=30'd256519562;
array2[12401]=30'd228216193;
array2[12402]=30'd231362949;
array2[12403]=30'd228216193;
array2[12404]=30'd231362949;
array2[12405]=30'd228216193;
array2[12406]=30'd228216193;
array2[12407]=30'd228216193;
array2[12408]=30'd228216193;
array2[12409]=30'd234504581;
array2[12410]=30'd231362949;
array2[12411]=30'd208120309;
array2[12412]=30'd768729747;
array2[12413]=30'd805398138;
array2[12414]=30'd819020415;
array2[12415]=30'd805398138;
array2[12416]=30'd805398138;
array2[12417]=30'd727851632;
array2[12418]=30'd190356956;
array2[12419]=30'd230307208;
array2[12420]=30'd234504581;
array2[12421]=30'd231362949;
array2[12422]=30'd256519562;
array2[12423]=30'd256519562;
array2[12424]=30'd228216193;
array2[12425]=30'd231362949;
array2[12426]=30'd231362949;
array2[12427]=30'd234504581;
array2[12428]=30'd228216193;
array2[12429]=30'd228216193;
array2[12430]=30'd227165569;
array2[12431]=30'd256519562;
array2[12432]=30'd472496545;
array2[12433]=30'd256519562;
array2[12434]=30'd231362949;
array2[12435]=30'd231364996;
array2[12436]=30'd231364996;
array2[12437]=30'd231362949;
array2[12438]=30'd212454818;
array2[12439]=30'd195647926;
array2[12440]=30'd179916222;
array2[12441]=30'd383147560;
array2[12442]=30'd672348794;
array2[12443]=30'd768729747;
array2[12444]=30'd819020415;
array2[12445]=30'd828452495;
array2[12446]=30'd828452495;
array2[12447]=30'd828452495;
array2[12448]=30'd851505800;
array2[12449]=30'd799112870;
array2[12450]=30'd727851632;
array2[12451]=30'd768729747;
array2[12452]=30'd770812573;
array2[12453]=30'd828452495;
array2[12454]=30'd828452495;
array2[12455]=30'd828452495;
array2[12456]=30'd819020415;
array2[12457]=30'd646130287;
array2[12458]=30'd506770009;
array2[12459]=30'd260631016;
array2[12460]=30'd257539480;
array2[12461]=30'd262793620;
array2[12462]=30'd262793620;
array2[12463]=30'd262793620;
array2[12464]=30'd238691720;
array2[12465]=30'd238691720;
array2[12466]=30'd228216193;
array2[12467]=30'd231362949;
array2[12468]=30'd229266819;
array2[12469]=30'd229266819;
array2[12470]=30'd231362949;
array2[12471]=30'd229266819;
array2[12472]=30'd231364996;
array2[12473]=30'd231362949;
array2[12474]=30'd231362949;
array2[12475]=30'd231362949;
array2[12476]=30'd231362949;
array2[12477]=30'd231362949;
array2[12478]=30'd231362949;
array2[12479]=30'd231362949;
array2[12480]=30'd193577377;
array2[12481]=30'd238691720;
array2[12482]=30'd238691720;
array2[12483]=30'd231362949;
array2[12484]=30'd232392085;
array2[12485]=30'd232392085;
array2[12486]=30'd232392085;
array2[12487]=30'd227159434;
array2[12488]=30'd232392085;
array2[12489]=30'd232392085;
array2[12490]=30'd232392085;
array2[12491]=30'd234499470;
array2[12492]=30'd232392085;
array2[12493]=30'd234499470;
array2[12494]=30'd232392085;
array2[12495]=30'd401193372;
array2[12496]=30'd405404052;
array2[12497]=30'd232392085;
array2[12498]=30'd238691720;
array2[12499]=30'd227159434;
array2[12500]=30'd238691720;
array2[12501]=30'd238691720;
array2[12502]=30'd234504581;
array2[12503]=30'd234499470;
array2[12504]=30'd238691720;
array2[12505]=30'd238691720;
array2[12506]=30'd231362949;
array2[12507]=30'd124307934;
array2[12508]=30'd450208341;
array2[12509]=30'd483727963;
array2[12510]=30'd483727963;
array2[12511]=30'd506770009;
array2[12512]=30'd762499681;
array2[12513]=30'd727851632;
array2[12514]=30'd190356956;
array2[12515]=30'd248105365;
array2[12516]=30'd232392085;
array2[12517]=30'd232392085;
array2[12518]=30'd338288022;
array2[12519]=30'd405404052;
array2[12520]=30'd262793620;
array2[12521]=30'd234504581;
array2[12522]=30'd234499470;
array2[12523]=30'd238691720;
array2[12524]=30'd238691720;
array2[12525]=30'd227159434;
array2[12526]=30'd238691720;
array2[12527]=30'd238691720;
array2[12528]=30'd256519562;
array2[12529]=30'd231364996;
array2[12530]=30'd229270912;
array2[12531]=30'd231364996;
array2[12532]=30'd231362949;
array2[12533]=30'd231362949;
array2[12534]=30'd231362949;
array2[12535]=30'd193577377;
array2[12536]=30'd179916222;
array2[12537]=30'd159912438;
array2[12538]=30'd407216718;
array2[12539]=30'd560184961;
array2[12540]=30'd678602388;
array2[12541]=30'd828452495;
array2[12542]=30'd851505800;
array2[12543]=30'd851505800;
array2[12544]=30'd851505800;
array2[12545]=30'd851505800;
array2[12546]=30'd858839683;
array2[12547]=30'd828452495;
array2[12548]=30'd858839683;
array2[12549]=30'd851505800;
array2[12550]=30'd851505800;
array2[12551]=30'd851505800;
array2[12552]=30'd851505800;
array2[12553]=30'd858839683;
array2[12554]=30'd770816666;
array2[12555]=30'd518272648;
array2[12556]=30'd260631016;
array2[12557]=30'd265928088;
array2[12558]=30'd262793620;
array2[12559]=30'd262793620;
array2[12560]=30'd238691720;
array2[12561]=30'd238691720;
array2[12562]=30'd227165569;
array2[12563]=30'd228216193;
array2[12564]=30'd229266819;
array2[12565]=30'd230317442;
array2[12566]=30'd231362949;
array2[12567]=30'd229266819;
array2[12568]=30'd231362949;
array2[12569]=30'd231362949;
array2[12570]=30'd229266819;
array2[12571]=30'd229266819;
array2[12572]=30'd231359873;
array2[12573]=30'd231362949;
array2[12574]=30'd231362949;
array2[12575]=30'd231362949;
array2[12576]=30'd307771998;
array2[12577]=30'd328674981;
array2[12578]=30'd307771998;
array2[12579]=30'd284737060;
array2[12580]=30'd357996288;
array2[12581]=30'd451191548;
array2[12582]=30'd451191548;
array2[12583]=30'd451191548;
array2[12584]=30'd451191548;
array2[12585]=30'd451191548;
array2[12586]=30'd451191548;
array2[12587]=30'd451191548;
array2[12588]=30'd451191548;
array2[12589]=30'd451191548;
array2[12590]=30'd461700935;
array2[12591]=30'd357996288;
array2[12592]=30'd302506616;
array2[12593]=30'd328674981;
array2[12594]=30'd302506616;
array2[12595]=30'd302506616;
array2[12596]=30'd328674981;
array2[12597]=30'd328674981;
array2[12598]=30'd302506616;
array2[12599]=30'd328674981;
array2[12600]=30'd302506616;
array2[12601]=30'd302506616;
array2[12602]=30'd284737060;
array2[12603]=30'd328674981;
array2[12604]=30'd357996288;
array2[12605]=30'd357996288;
array2[12606]=30'd357996288;
array2[12607]=30'd287786593;
array2[12608]=30'd483727963;
array2[12609]=30'd481587821;
array2[12610]=30'd287786593;
array2[12611]=30'd357996288;
array2[12612]=30'd395649781;
array2[12613]=30'd390446940;
array2[12614]=30'd395649781;
array2[12615]=30'd328674981;
array2[12616]=30'd328674981;
array2[12617]=30'd328674981;
array2[12618]=30'd302506616;
array2[12619]=30'd302506616;
array2[12620]=30'd302506616;
array2[12621]=30'd302506616;
array2[12622]=30'd302506616;
array2[12623]=30'd307771998;
array2[12624]=30'd280568333;
array2[12625]=30'd227159434;
array2[12626]=30'd179916222;
array2[12627]=30'd179916222;
array2[12628]=30'd179916222;
array2[12629]=30'd179916222;
array2[12630]=30'd179916222;
array2[12631]=30'd407216718;
array2[12632]=30'd560184961;
array2[12633]=30'd606320275;
array2[12634]=30'd631447172;
array2[12635]=30'd631447172;
array2[12636]=30'd560184961;
array2[12637]=30'd560184961;
array2[12638]=30'd646130287;
array2[12639]=30'd768729747;
array2[12640]=30'd828452495;
array2[12641]=30'd858839683;
array2[12642]=30'd851505800;
array2[12643]=30'd858839683;
array2[12644]=30'd851505800;
array2[12645]=30'd851505800;
array2[12646]=30'd828452495;
array2[12647]=30'd851505800;
array2[12648]=30'd858839683;
array2[12649]=30'd858839683;
array2[12650]=30'd851505800;
array2[12651]=30'd770816666;
array2[12652]=30'd518272648;
array2[12653]=30'd193577377;
array2[12654]=30'd238691720;
array2[12655]=30'd262793620;
array2[12656]=30'd238691720;
array2[12657]=30'd238691720;
array2[12658]=30'd238691720;
array2[12659]=30'd227165569;
array2[12660]=30'd231362949;
array2[12661]=30'd231362949;
array2[12662]=30'd231362949;
array2[12663]=30'd230317442;
array2[12664]=30'd229266819;
array2[12665]=30'd229266819;
array2[12666]=30'd231362949;
array2[12667]=30'd231362949;
array2[12668]=30'd231362949;
array2[12669]=30'd231362949;
array2[12670]=30'd231362949;
array2[12671]=30'd231362949;
array2[12672]=30'd390446940;
array2[12673]=30'd429185963;
array2[12674]=30'd429185963;
array2[12675]=30'd409311115;
array2[12676]=30'd429185963;
array2[12677]=30'd429185963;
array2[12678]=30'd409311115;
array2[12679]=30'd429185963;
array2[12680]=30'd429185963;
array2[12681]=30'd429185963;
array2[12682]=30'd429185963;
array2[12683]=30'd409311115;
array2[12684]=30'd429185963;
array2[12685]=30'd429185963;
array2[12686]=30'd429185963;
array2[12687]=30'd409311115;
array2[12688]=30'd429185963;
array2[12689]=30'd409311115;
array2[12690]=30'd409311115;
array2[12691]=30'd409311115;
array2[12692]=30'd409311115;
array2[12693]=30'd409311115;
array2[12694]=30'd409311115;
array2[12695]=30'd409311115;
array2[12696]=30'd429185963;
array2[12697]=30'd409311115;
array2[12698]=30'd409311115;
array2[12699]=30'd429185963;
array2[12700]=30'd429185963;
array2[12701]=30'd429185963;
array2[12702]=30'd429185963;
array2[12703]=30'd328674981;
array2[12704]=30'd338018898;
array2[12705]=30'd357913199;
array2[12706]=30'd287786593;
array2[12707]=30'd461700935;
array2[12708]=30'd409311115;
array2[12709]=30'd409311115;
array2[12710]=30'd429185963;
array2[12711]=30'd409311115;
array2[12712]=30'd409311115;
array2[12713]=30'd409311115;
array2[12714]=30'd409311115;
array2[12715]=30'd409311115;
array2[12716]=30'd409311115;
array2[12717]=30'd409311115;
array2[12718]=30'd409311115;
array2[12719]=30'd357996288;
array2[12720]=30'd218607140;
array2[12721]=30'd249001484;
array2[12722]=30'd631447172;
array2[12723]=30'd677571193;
array2[12724]=30'd331763301;
array2[12725]=30'd331763301;
array2[12726]=30'd331763301;
array2[12727]=30'd606320275;
array2[12728]=30'd732038833;
array2[12729]=30'd770812573;
array2[12730]=30'd770812573;
array2[12731]=30'd732038833;
array2[12732]=30'd732038833;
array2[12733]=30'd713179821;
array2[12734]=30'd604201637;
array2[12735]=30'd565444213;
array2[12736]=30'd646130287;
array2[12737]=30'd851505800;
array2[12738]=30'd851505800;
array2[12739]=30'd851505800;
array2[12740]=30'd851505800;
array2[12741]=30'd858839683;
array2[12742]=30'd851505800;
array2[12743]=30'd851505800;
array2[12744]=30'd858839683;
array2[12745]=30'd858839683;
array2[12746]=30'd858839683;
array2[12747]=30'd851505800;
array2[12748]=30'd727851632;
array2[12749]=30'd179916222;
array2[12750]=30'd227159434;
array2[12751]=30'd262793620;
array2[12752]=30'd262793620;
array2[12753]=30'd227159434;
array2[12754]=30'd234504581;
array2[12755]=30'd228216193;
array2[12756]=30'd231364996;
array2[12757]=30'd231364996;
array2[12758]=30'd228216193;
array2[12759]=30'd231362949;
array2[12760]=30'd230317442;
array2[12761]=30'd231362949;
array2[12762]=30'd230317442;
array2[12763]=30'd229266819;
array2[12764]=30'd231362949;
array2[12765]=30'd231362949;
array2[12766]=30'd234504581;
array2[12767]=30'd231362949;
array2[12768]=30'd461700935;
array2[12769]=30'd423950257;
array2[12770]=30'd423950257;
array2[12771]=30'd423950257;
array2[12772]=30'd423950257;
array2[12773]=30'd426044336;
array2[12774]=30'd423950257;
array2[12775]=30'd423950257;
array2[12776]=30'd423950257;
array2[12777]=30'd423950257;
array2[12778]=30'd426044336;
array2[12779]=30'd423950257;
array2[12780]=30'd426044336;
array2[12781]=30'd423950257;
array2[12782]=30'd423950257;
array2[12783]=30'd423950257;
array2[12784]=30'd426044336;
array2[12785]=30'd423950257;
array2[12786]=30'd423950257;
array2[12787]=30'd423950257;
array2[12788]=30'd423950257;
array2[12789]=30'd423950257;
array2[12790]=30'd426044336;
array2[12791]=30'd423950257;
array2[12792]=30'd423950257;
array2[12793]=30'd423950257;
array2[12794]=30'd426044336;
array2[12795]=30'd426044336;
array2[12796]=30'd423950257;
array2[12797]=30'd426044336;
array2[12798]=30'd429185963;
array2[12799]=30'd328674981;
array2[12800]=30'd338018898;
array2[12801]=30'd331763301;
array2[12802]=30'd218607140;
array2[12803]=30'd218607140;
array2[12804]=30'd218607140;
array2[12805]=30'd218607140;
array2[12806]=30'd461700935;
array2[12807]=30'd423950257;
array2[12808]=30'd423950257;
array2[12809]=30'd423950257;
array2[12810]=30'd423950257;
array2[12811]=30'd426044336;
array2[12812]=30'd429185963;
array2[12813]=30'd390446940;
array2[12814]=30'd299264555;
array2[12815]=30'd295074390;
array2[12816]=30'd560184961;
array2[12817]=30'd770812573;
array2[12818]=30'd828452495;
array2[12819]=30'd768729747;
array2[12820]=30'd434416250;
array2[12821]=30'd375721588;
array2[12822]=30'd375721588;
array2[12823]=30'd677571193;
array2[12824]=30'd828452495;
array2[12825]=30'd851505800;
array2[12826]=30'd851505800;
array2[12827]=30'd851505800;
array2[12828]=30'd851505800;
array2[12829]=30'd858839683;
array2[12830]=30'd858839683;
array2[12831]=30'd828452495;
array2[12832]=30'd828452495;
array2[12833]=30'd851505800;
array2[12834]=30'd858839683;
array2[12835]=30'd858839683;
array2[12836]=30'd851505800;
array2[12837]=30'd858839683;
array2[12838]=30'd858839683;
array2[12839]=30'd865130113;
array2[12840]=30'd858839683;
array2[12841]=30'd851505800;
array2[12842]=30'd805398138;
array2[12843]=30'd805398138;
array2[12844]=30'd828452495;
array2[12845]=30'd483727963;
array2[12846]=30'd207191473;
array2[12847]=30'd262793620;
array2[12848]=30'd262793620;
array2[12849]=30'd238691720;
array2[12850]=30'd238691720;
array2[12851]=30'd228216193;
array2[12852]=30'd230317442;
array2[12853]=30'd231364996;
array2[12854]=30'd231364996;
array2[12855]=30'd231362949;
array2[12856]=30'd231362949;
array2[12857]=30'd228216193;
array2[12858]=30'd229266819;
array2[12859]=30'd229266819;
array2[12860]=30'd231359873;
array2[12861]=30'd231359873;
array2[12862]=30'd234504581;
array2[12863]=30'd231362949;
array2[12864]=30'd461700935;
array2[12865]=30'd493111164;
array2[12866]=30'd493111164;
array2[12867]=30'd435467177;
array2[12868]=30'd582196031;
array2[12869]=30'd582196031;
array2[12870]=30'd582196031;
array2[12871]=30'd582196031;
array2[12872]=30'd635645720;
array2[12873]=30'd582196031;
array2[12874]=30'd582196031;
array2[12875]=30'd635645720;
array2[12876]=30'd582196031;
array2[12877]=30'd635645720;
array2[12878]=30'd672324351;
array2[12879]=30'd582196031;
array2[12880]=30'd493111164;
array2[12881]=30'd493111164;
array2[12882]=30'd493111164;
array2[12883]=30'd493111164;
array2[12884]=30'd493111164;
array2[12885]=30'd493111164;
array2[12886]=30'd493111164;
array2[12887]=30'd493111164;
array2[12888]=30'd493111164;
array2[12889]=30'd493111164;
array2[12890]=30'd435467177;
array2[12891]=30'd582196031;
array2[12892]=30'd582196031;
array2[12893]=30'd582196031;
array2[12894]=30'd635645720;
array2[12895]=30'd339090072;
array2[12896]=30'd265736724;
array2[12897]=30'd295074390;
array2[12898]=30'd295074390;
array2[12899]=30'd338018898;
array2[12900]=30'd357913199;
array2[12901]=30'd222764576;
array2[12902]=30'd558174979;
array2[12903]=30'd493111164;
array2[12904]=30'd493111164;
array2[12905]=30'd493111164;
array2[12906]=30'd493111164;
array2[12907]=30'd493111164;
array2[12908]=30'd390446940;
array2[12909]=30'd295074390;
array2[12910]=30'd331763301;
array2[12911]=30'd357913199;
array2[12912]=30'd672348794;
array2[12913]=30'd851505800;
array2[12914]=30'd851505800;
array2[12915]=30'd805398138;
array2[12916]=30'd518272648;
array2[12917]=30'd375721588;
array2[12918]=30'd375721588;
array2[12919]=30'd727851632;
array2[12920]=30'd858839683;
array2[12921]=30'd851505800;
array2[12922]=30'd858839683;
array2[12923]=30'd851505800;
array2[12924]=30'd851505800;
array2[12925]=30'd851505800;
array2[12926]=30'd858839683;
array2[12927]=30'd858839683;
array2[12928]=30'd858839683;
array2[12929]=30'd851505800;
array2[12930]=30'd865130113;
array2[12931]=30'd865130113;
array2[12932]=30'd858839683;
array2[12933]=30'd858839683;
array2[12934]=30'd851505800;
array2[12935]=30'd858839683;
array2[12936]=30'd865130113;
array2[12937]=30'd819020415;
array2[12938]=30'd401997362;
array2[12939]=30'd401997362;
array2[12940]=30'd819020415;
array2[12941]=30'd566515308;
array2[12942]=30'd207191473;
array2[12943]=30'd271165847;
array2[12944]=30'd265928088;
array2[12945]=30'd265928088;
array2[12946]=30'd234504581;
array2[12947]=30'd234504581;
array2[12948]=30'd228216193;
array2[12949]=30'd231362949;
array2[12950]=30'd230317442;
array2[12951]=30'd234504581;
array2[12952]=30'd231364996;
array2[12953]=30'd229266819;
array2[12954]=30'd229266819;
array2[12955]=30'd231362949;
array2[12956]=30'd231362949;
array2[12957]=30'd231362949;
array2[12958]=30'd231362949;
array2[12959]=30'd231362949;
array2[12960]=30'd601041592;
array2[12961]=30'd672324351;
array2[12962]=30'd718417640;
array2[12963]=30'd672324351;
array2[12964]=30'd718417640;
array2[12965]=30'd718417640;
array2[12966]=30'd718417640;
array2[12967]=30'd718417640;
array2[12968]=30'd718417640;
array2[12969]=30'd718417640;
array2[12970]=30'd718417640;
array2[12971]=30'd728897252;
array2[12972]=30'd728897252;
array2[12973]=30'd718417640;
array2[12974]=30'd728897252;
array2[12975]=30'd718417640;
array2[12976]=30'd672324351;
array2[12977]=30'd672324351;
array2[12978]=30'd718417640;
array2[12979]=30'd718417640;
array2[12980]=30'd672324351;
array2[12981]=30'd718417640;
array2[12982]=30'd718417640;
array2[12983]=30'd672324351;
array2[12984]=30'd718417640;
array2[12985]=30'd672324351;
array2[12986]=30'd672324351;
array2[12987]=30'd718417640;
array2[12988]=30'd728897252;
array2[12989]=30'd718417640;
array2[12990]=30'd718417640;
array2[12991]=30'd539218630;
array2[12992]=30'd481587821;
array2[12993]=30'd481587821;
array2[12994]=30'd481587821;
array2[12995]=30'd450208341;
array2[12996]=30'd331763301;
array2[12997]=30'd299264555;
array2[12998]=30'd646169309;
array2[12999]=30'd672324351;
array2[13000]=30'd718417640;
array2[13001]=30'd718417640;
array2[13002]=30'd672324351;
array2[13003]=30'd601041592;
array2[13004]=30'd449120871;
array2[13005]=30'd357913199;
array2[13006]=30'd375721588;
array2[13007]=30'd375721588;
array2[13008]=30'd646130287;
array2[13009]=30'd858839683;
array2[13010]=30'd851505800;
array2[13011]=30'd851505800;
array2[13012]=30'd711090860;
array2[13013]=30'd450208341;
array2[13014]=30'd375721588;
array2[13015]=30'd727851632;
array2[13016]=30'd828452495;
array2[13017]=30'd851505800;
array2[13018]=30'd858839683;
array2[13019]=30'd858839683;
array2[13020]=30'd858839683;
array2[13021]=30'd858839683;
array2[13022]=30'd865130113;
array2[13023]=30'd865130113;
array2[13024]=30'd865130113;
array2[13025]=30'd858839683;
array2[13026]=30'd858839683;
array2[13027]=30'd858839683;
array2[13028]=30'd851505800;
array2[13029]=30'd865130113;
array2[13030]=30'd858839683;
array2[13031]=30'd865130113;
array2[13032]=30'd858839683;
array2[13033]=30'd819020415;
array2[13034]=30'd401997362;
array2[13035]=30'd383147560;
array2[13036]=30'd823228019;
array2[13037]=30'd566515308;
array2[13038]=30'd207191473;
array2[13039]=30'd265928088;
array2[13040]=30'd262793620;
array2[13041]=30'd262793620;
array2[13042]=30'd234504581;
array2[13043]=30'd227165569;
array2[13044]=30'd234504581;
array2[13045]=30'd231362949;
array2[13046]=30'd231362949;
array2[13047]=30'd227165569;
array2[13048]=30'd231362949;
array2[13049]=30'd229270912;
array2[13050]=30'd230317442;
array2[13051]=30'd231362949;
array2[13052]=30'd228216193;
array2[13053]=30'd229266819;
array2[13054]=30'd229266819;
array2[13055]=30'd231362949;
array2[13056]=30'd678602388;
array2[13057]=30'd728897252;
array2[13058]=30'd728897252;
array2[13059]=30'd728897252;
array2[13060]=30'd728897252;
array2[13061]=30'd728897252;
array2[13062]=30'd728897252;
array2[13063]=30'd728897252;
array2[13064]=30'd728897252;
array2[13065]=30'd728897252;
array2[13066]=30'd728897252;
array2[13067]=30'd728897252;
array2[13068]=30'd728897252;
array2[13069]=30'd728897252;
array2[13070]=30'd728897252;
array2[13071]=30'd728897252;
array2[13072]=30'd728897252;
array2[13073]=30'd728897252;
array2[13074]=30'd728897252;
array2[13075]=30'd728897252;
array2[13076]=30'd728897252;
array2[13077]=30'd728897252;
array2[13078]=30'd728897252;
array2[13079]=30'd728897252;
array2[13080]=30'd728897252;
array2[13081]=30'd728897252;
array2[13082]=30'd728897252;
array2[13083]=30'd728897252;
array2[13084]=30'd728897252;
array2[13085]=30'd728897252;
array2[13086]=30'd728897252;
array2[13087]=30'd728897252;
array2[13088]=30'd728897252;
array2[13089]=30'd728897252;
array2[13090]=30'd728897252;
array2[13091]=30'd601041592;
array2[13092]=30'd299264555;
array2[13093]=30'd299264555;
array2[13094]=30'd646169309;
array2[13095]=30'd718417640;
array2[13096]=30'd718417640;
array2[13097]=30'd718417640;
array2[13098]=30'd601041592;
array2[13099]=30'd518272648;
array2[13100]=30'd713179821;
array2[13101]=30'd631447172;
array2[13102]=30'd375721588;
array2[13103]=30'd375721588;
array2[13104]=30'd631447172;
array2[13105]=30'd828452495;
array2[13106]=30'd858839683;
array2[13107]=30'd858839683;
array2[13108]=30'd819020415;
array2[13109]=30'd606320275;
array2[13110]=30'd375721588;
array2[13111]=30'd678602388;
array2[13112]=30'd819020415;
array2[13113]=30'd858839683;
array2[13114]=30'd851505800;
array2[13115]=30'd858839683;
array2[13116]=30'd851505800;
array2[13117]=30'd865130113;
array2[13118]=30'd858839683;
array2[13119]=30'd858839683;
array2[13120]=30'd858839683;
array2[13121]=30'd858839683;
array2[13122]=30'd851505800;
array2[13123]=30'd858839683;
array2[13124]=30'd851505800;
array2[13125]=30'd865130113;
array2[13126]=30'd865130113;
array2[13127]=30'd851505800;
array2[13128]=30'd858839683;
array2[13129]=30'd819020415;
array2[13130]=30'd450208341;
array2[13131]=30'd401997362;
array2[13132]=30'd805398138;
array2[13133]=30'd566515308;
array2[13134]=30'd195647926;
array2[13135]=30'd265928088;
array2[13136]=30'd232392085;
array2[13137]=30'd262793620;
array2[13138]=30'd262793620;
array2[13139]=30'd227165569;
array2[13140]=30'd238691720;
array2[13141]=30'd228216193;
array2[13142]=30'd231362949;
array2[13143]=30'd231362949;
array2[13144]=30'd230317442;
array2[13145]=30'd230317442;
array2[13146]=30'd229270912;
array2[13147]=30'd231362949;
array2[13148]=30'd231362949;
array2[13149]=30'd228216193;
array2[13150]=30'd229266819;
array2[13151]=30'd229266819;
array2[13152]=30'd678602388;
array2[13153]=30'd758240964;
array2[13154]=30'd758240964;
array2[13155]=30'd758240964;
array2[13156]=30'd799112870;
array2[13157]=30'd828452495;
array2[13158]=30'd828452495;
array2[13159]=30'd828452495;
array2[13160]=30'd828452495;
array2[13161]=30'd828452495;
array2[13162]=30'd828452495;
array2[13163]=30'd828452495;
array2[13164]=30'd828452495;
array2[13165]=30'd828452495;
array2[13166]=30'd851505800;
array2[13167]=30'd828452495;
array2[13168]=30'd758240964;
array2[13169]=30'd799112870;
array2[13170]=30'd758240964;
array2[13171]=30'd758240964;
array2[13172]=30'd758240964;
array2[13173]=30'd799112870;
array2[13174]=30'd758240964;
array2[13175]=30'd758240964;
array2[13176]=30'd758240964;
array2[13177]=30'd758240964;
array2[13178]=30'd728897252;
array2[13179]=30'd758240964;
array2[13180]=30'd828452495;
array2[13181]=30'd828452495;
array2[13182]=30'd828452495;
array2[13183]=30'd828452495;
array2[13184]=30'd828452495;
array2[13185]=30'd828452495;
array2[13186]=30'd828452495;
array2[13187]=30'd727851632;
array2[13188]=30'd299264555;
array2[13189]=30'd295074390;
array2[13190]=30'd338018898;
array2[13191]=30'd407216718;
array2[13192]=30'd407216718;
array2[13193]=30'd375721588;
array2[13194]=30'd481587821;
array2[13195]=30'd768729747;
array2[13196]=30'd828452495;
array2[13197]=30'd819020415;
array2[13198]=30'd606320275;
array2[13199]=30'd375721588;
array2[13200]=30'd434416250;
array2[13201]=30'd727851632;
array2[13202]=30'd858839683;
array2[13203]=30'd851505800;
array2[13204]=30'd851505800;
array2[13205]=30'd713179821;
array2[13206]=30'd434416250;
array2[13207]=30'd764529268;
array2[13208]=30'd828452495;
array2[13209]=30'd851505800;
array2[13210]=30'd851505800;
array2[13211]=30'd858839683;
array2[13212]=30'd858839683;
array2[13213]=30'd858839683;
array2[13214]=30'd858839683;
array2[13215]=30'd865130113;
array2[13216]=30'd858839683;
array2[13217]=30'd865130113;
array2[13218]=30'd858839683;
array2[13219]=30'd858839683;
array2[13220]=30'd851505800;
array2[13221]=30'd770812573;
array2[13222]=30'd646169309;
array2[13223]=30'd732038833;
array2[13224]=30'd828452495;
array2[13225]=30'd819020415;
array2[13226]=30'd485780117;
array2[13227]=30'd560184961;
array2[13228]=30'd799112870;
array2[13229]=30'd711090860;
array2[13230]=30'd444954173;
array2[13231]=30'd190356956;
array2[13232]=30'd228181405;
array2[13233]=30'd262793620;
array2[13234]=30'd262793620;
array2[13235]=30'd234504581;
array2[13236]=30'd234504581;
array2[13237]=30'd231362949;
array2[13238]=30'd231362949;
array2[13239]=30'd231364996;
array2[13240]=30'd228216193;
array2[13241]=30'd229266819;
array2[13242]=30'd231362949;
array2[13243]=30'd231364996;
array2[13244]=30'd229266819;
array2[13245]=30'd229266819;
array2[13246]=30'd231362949;
array2[13247]=30'd234504581;
array2[13248]=30'd762499681;
array2[13249]=30'd865130113;
array2[13250]=30'd865130113;
array2[13251]=30'd865130113;
array2[13252]=30'd906004072;
array2[13253]=30'd906004072;
array2[13254]=30'd906004072;
array2[13255]=30'd906004072;
array2[13256]=30'd906004072;
array2[13257]=30'd906004072;
array2[13258]=30'd906004072;
array2[13259]=30'd906004072;
array2[13260]=30'd906004072;
array2[13261]=30'd906004072;
array2[13262]=30'd906004072;
array2[13263]=30'd906004072;
array2[13264]=30'd906004072;
array2[13265]=30'd906004072;
array2[13266]=30'd906004072;
array2[13267]=30'd865130113;
array2[13268]=30'd865130113;
array2[13269]=30'd906004072;
array2[13270]=30'd865130113;
array2[13271]=30'd865130113;
array2[13272]=30'd865130113;
array2[13273]=30'd865130113;
array2[13274]=30'd865130113;
array2[13275]=30'd906004072;
array2[13276]=30'd906004072;
array2[13277]=30'd906004072;
array2[13278]=30'd906004072;
array2[13279]=30'd906004072;
array2[13280]=30'd906004072;
array2[13281]=30'd906004072;
array2[13282]=30'd906004072;
array2[13283]=30'd749877860;
array2[13284]=30'd347490866;
array2[13285]=30'd347490866;
array2[13286]=30'd347490866;
array2[13287]=30'd347490866;
array2[13288]=30'd319215128;
array2[13289]=30'd449120871;
array2[13290]=30'd764529268;
array2[13291]=30'd828452495;
array2[13292]=30'd851505800;
array2[13293]=30'd851505800;
array2[13294]=30'd770812573;
array2[13295]=30'd606320275;
array2[13296]=30'd449120871;
array2[13297]=30'd727851632;
array2[13298]=30'd851505800;
array2[13299]=30'd851505800;
array2[13300]=30'd851505800;
array2[13301]=30'd828452495;
array2[13302]=30'd805398138;
array2[13303]=30'd819020415;
array2[13304]=30'd858839683;
array2[13305]=30'd851505800;
array2[13306]=30'd851505800;
array2[13307]=30'd851505800;
array2[13308]=30'd865130113;
array2[13309]=30'd858839683;
array2[13310]=30'd865130113;
array2[13311]=30'd858839683;
array2[13312]=30'd858839683;
array2[13313]=30'd858839683;
array2[13314]=30'd865130113;
array2[13315]=30'd858839683;
array2[13316]=30'd770816666;
array2[13317]=30'd539218630;
array2[13318]=30'd409311115;
array2[13319]=30'd558174979;
array2[13320]=30'd732038833;
array2[13321]=30'd828452495;
array2[13322]=30'd768729747;
array2[13323]=30'd770812573;
array2[13324]=30'd851505800;
array2[13325]=30'd828452495;
array2[13326]=30'd764529268;
array2[13327]=30'd319215128;
array2[13328]=30'd228181405;
array2[13329]=30'd262793620;
array2[13330]=30'd227159434;
array2[13331]=30'd227165569;
array2[13332]=30'd231362949;
array2[13333]=30'd229266819;
array2[13334]=30'd234504581;
array2[13335]=30'd231364996;
array2[13336]=30'd229266819;
array2[13337]=30'd229266819;
array2[13338]=30'd231362949;
array2[13339]=30'd231362949;
array2[13340]=30'd231362949;
array2[13341]=30'd229266819;
array2[13342]=30'd231362949;
array2[13343]=30'd229266819;
array2[13344]=30'd764529268;
array2[13345]=30'd906004072;
array2[13346]=30'd906004072;
array2[13347]=30'd906004072;
array2[13348]=30'd906004072;
array2[13349]=30'd906004072;
array2[13350]=30'd906004072;
array2[13351]=30'd906004072;
array2[13352]=30'd906004072;
array2[13353]=30'd906004072;
array2[13354]=30'd906004072;
array2[13355]=30'd906004072;
array2[13356]=30'd906004072;
array2[13357]=30'd906004072;
array2[13358]=30'd906004072;
array2[13359]=30'd906004072;
array2[13360]=30'd906004072;
array2[13361]=30'd906004072;
array2[13362]=30'd906004072;
array2[13363]=30'd906004072;
array2[13364]=30'd906004072;
array2[13365]=30'd906004072;
array2[13366]=30'd906004072;
array2[13367]=30'd906004072;
array2[13368]=30'd906004072;
array2[13369]=30'd906004072;
array2[13370]=30'd906004072;
array2[13371]=30'd906004072;
array2[13372]=30'd906004072;
array2[13373]=30'd906004072;
array2[13374]=30'd906004072;
array2[13375]=30'd906004072;
array2[13376]=30'd906004072;
array2[13377]=30'd906004072;
array2[13378]=30'd906004072;
array2[13379]=30'd906004072;
array2[13380]=30'd823228019;
array2[13381]=30'd823228019;
array2[13382]=30'd823228019;
array2[13383]=30'd823228019;
array2[13384]=30'd678604396;
array2[13385]=30'd506770009;
array2[13386]=30'd858839683;
array2[13387]=30'd851505800;
array2[13388]=30'd851505800;
array2[13389]=30'd858839683;
array2[13390]=30'd858839683;
array2[13391]=30'd828452495;
array2[13392]=30'd819020415;
array2[13393]=30'd851505800;
array2[13394]=30'd851505800;
array2[13395]=30'd851505800;
array2[13396]=30'd858839683;
array2[13397]=30'd858839683;
array2[13398]=30'd858839683;
array2[13399]=30'd865130113;
array2[13400]=30'd858839683;
array2[13401]=30'd851505800;
array2[13402]=30'd858839683;
array2[13403]=30'd851505800;
array2[13404]=30'd865130113;
array2[13405]=30'd858839683;
array2[13406]=30'd858839683;
array2[13407]=30'd858839683;
array2[13408]=30'd858839683;
array2[13409]=30'd865130113;
array2[13410]=30'd858839683;
array2[13411]=30'd851505800;
array2[13412]=30'd451191548;
array2[13413]=30'd395649781;
array2[13414]=30'd451191548;
array2[13415]=30'd409311115;
array2[13416]=30'd558174979;
array2[13417]=30'd770812573;
array2[13418]=30'd851505800;
array2[13419]=30'd828452495;
array2[13420]=30'd851505800;
array2[13421]=30'd858839683;
array2[13422]=30'd828452495;
array2[13423]=30'd347490866;
array2[13424]=30'd212454818;
array2[13425]=30'd262793620;
array2[13426]=30'd227165569;
array2[13427]=30'd228216193;
array2[13428]=30'd228216193;
array2[13429]=30'd231362949;
array2[13430]=30'd231362949;
array2[13431]=30'd231364996;
array2[13432]=30'd231364996;
array2[13433]=30'd231362949;
array2[13434]=30'd228216193;
array2[13435]=30'd228216193;
array2[13436]=30'd230317442;
array2[13437]=30'd231362949;
array2[13438]=30'd231359873;
array2[13439]=30'd231362949;
array2[13440]=30'd729975381;
array2[13441]=30'd832648722;
array2[13442]=30'd832648722;
array2[13443]=30'd906004072;
array2[13444]=30'd783393281;
array2[13445]=30'd736232864;
array2[13446]=30'd736232864;
array2[13447]=30'd736232864;
array2[13448]=30'd736232864;
array2[13449]=30'd736232864;
array2[13450]=30'd736232864;
array2[13451]=30'd736232864;
array2[13452]=30'd736232864;
array2[13453]=30'd736232864;
array2[13454]=30'd736232864;
array2[13455]=30'd783393281;
array2[13456]=30'd832648722;
array2[13457]=30'd832648722;
array2[13458]=30'd832648722;
array2[13459]=30'd832648722;
array2[13460]=30'd832648722;
array2[13461]=30'd832648722;
array2[13462]=30'd832648722;
array2[13463]=30'd832648722;
array2[13464]=30'd832648722;
array2[13465]=30'd832648722;
array2[13466]=30'd906004072;
array2[13467]=30'd815880708;
array2[13468]=30'd736232864;
array2[13469]=30'd736232864;
array2[13470]=30'd736232864;
array2[13471]=30'd736232864;
array2[13472]=30'd736232864;
array2[13473]=30'd736232864;
array2[13474]=30'd736232864;
array2[13475]=30'd736232864;
array2[13476]=30'd736232864;
array2[13477]=30'd736232864;
array2[13478]=30'd736232864;
array2[13479]=30'd783393281;
array2[13480]=30'd401997362;
array2[13481]=30'd819020415;
array2[13482]=30'd851505800;
array2[13483]=30'd865130113;
array2[13484]=30'd858839683;
array2[13485]=30'd851505800;
array2[13486]=30'd858839683;
array2[13487]=30'd851505800;
array2[13488]=30'd865130113;
array2[13489]=30'd865130113;
array2[13490]=30'd858839683;
array2[13491]=30'd858839683;
array2[13492]=30'd858839683;
array2[13493]=30'd858839683;
array2[13494]=30'd858839683;
array2[13495]=30'd865130113;
array2[13496]=30'd858839683;
array2[13497]=30'd858839683;
array2[13498]=30'd858839683;
array2[13499]=30'd865130113;
array2[13500]=30'd858839683;
array2[13501]=30'd858839683;
array2[13502]=30'd865130113;
array2[13503]=30'd858839683;
array2[13504]=30'd858839683;
array2[13505]=30'd865130113;
array2[13506]=30'd858839683;
array2[13507]=30'd858839683;
array2[13508]=30'd539218630;
array2[13509]=30'd395649781;
array2[13510]=30'd395649781;
array2[13511]=30'd451191548;
array2[13512]=30'd461700935;
array2[13513]=30'd770812573;
array2[13514]=30'd851505800;
array2[13515]=30'd851505800;
array2[13516]=30'd851505800;
array2[13517]=30'd819020415;
array2[13518]=30'd711090860;
array2[13519]=30'd299264555;
array2[13520]=30'd212454818;
array2[13521]=30'd238691720;
array2[13522]=30'd234504581;
array2[13523]=30'd229266819;
array2[13524]=30'd230317442;
array2[13525]=30'd231362949;
array2[13526]=30'd227165569;
array2[13527]=30'd231359873;
array2[13528]=30'd230317442;
array2[13529]=30'd231362949;
array2[13530]=30'd231362949;
array2[13531]=30'd231362949;
array2[13532]=30'd229270912;
array2[13533]=30'd231362949;
array2[13534]=30'd231359873;
array2[13535]=30'd231362949;
array2[13536]=30'd582318295;
array2[13537]=30'd690121052;
array2[13538]=30'd690121052;
array2[13539]=30'd690121052;
array2[13540]=30'd639824186;
array2[13541]=30'd637725975;
array2[13542]=30'd637725975;
array2[13543]=30'd637725975;
array2[13544]=30'd637725975;
array2[13545]=30'd637725975;
array2[13546]=30'd637725975;
array2[13547]=30'd637725975;
array2[13548]=30'd637725975;
array2[13549]=30'd637725975;
array2[13550]=30'd615715061;
array2[13551]=30'd637725975;
array2[13552]=30'd690121052;
array2[13553]=30'd690121052;
array2[13554]=30'd690121052;
array2[13555]=30'd690121052;
array2[13556]=30'd690121052;
array2[13557]=30'd690121052;
array2[13558]=30'd690121052;
array2[13559]=30'd690121052;
array2[13560]=30'd690121052;
array2[13561]=30'd690121052;
array2[13562]=30'd690121052;
array2[13563]=30'd690121052;
array2[13564]=30'd637725975;
array2[13565]=30'd637725975;
array2[13566]=30'd637725975;
array2[13567]=30'd637725975;
array2[13568]=30'd637725975;
array2[13569]=30'd637725975;
array2[13570]=30'd637725975;
array2[13571]=30'd637725975;
array2[13572]=30'd637725975;
array2[13573]=30'd615715061;
array2[13574]=30'd637725975;
array2[13575]=30'd639824186;
array2[13576]=30'd401997362;
array2[13577]=30'd858839683;
array2[13578]=30'd851505800;
array2[13579]=30'd851505800;
array2[13580]=30'd858839683;
array2[13581]=30'd858839683;
array2[13582]=30'd858839683;
array2[13583]=30'd858839683;
array2[13584]=30'd858839683;
array2[13585]=30'd865130113;
array2[13586]=30'd858839683;
array2[13587]=30'd858839683;
array2[13588]=30'd858839683;
array2[13589]=30'd865130113;
array2[13590]=30'd858839683;
array2[13591]=30'd858839683;
array2[13592]=30'd858839683;
array2[13593]=30'd858839683;
array2[13594]=30'd858839683;
array2[13595]=30'd858839683;
array2[13596]=30'd858839683;
array2[13597]=30'd858839683;
array2[13598]=30'd865130113;
array2[13599]=30'd858839683;
array2[13600]=30'd858839683;
array2[13601]=30'd865130113;
array2[13602]=30'd865130113;
array2[13603]=30'd858839683;
array2[13604]=30'd799112870;
array2[13605]=30'd601041592;
array2[13606]=30'd451191548;
array2[13607]=30'd537140990;
array2[13608]=30'd713179821;
array2[13609]=30'd828452495;
array2[13610]=30'd851505800;
array2[13611]=30'd851505800;
array2[13612]=30'd858839683;
array2[13613]=30'd711090860;
array2[13614]=30'd483727963;
array2[13615]=30'd179916222;
array2[13616]=30'd220861839;
array2[13617]=30'd227165569;
array2[13618]=30'd231362949;
array2[13619]=30'd231364996;
array2[13620]=30'd228216193;
array2[13621]=30'd231362949;
array2[13622]=30'd231364996;
array2[13623]=30'd231362949;
array2[13624]=30'd231362949;
array2[13625]=30'd231362949;
array2[13626]=30'd234504581;
array2[13627]=30'd231362949;
array2[13628]=30'd231364996;
array2[13629]=30'd228216193;
array2[13630]=30'd231362949;
array2[13631]=30'd231362949;
array2[13632]=30'd559300847;
array2[13633]=30'd611520752;
array2[13634]=30'd615715061;
array2[13635]=30'd611520752;
array2[13636]=30'd611520752;
array2[13637]=30'd611520752;
array2[13638]=30'd611520752;
array2[13639]=30'd615715061;
array2[13640]=30'd611520752;
array2[13641]=30'd611520752;
array2[13642]=30'd615715061;
array2[13643]=30'd611520752;
array2[13644]=30'd611520752;
array2[13645]=30'd615715061;
array2[13646]=30'd611520752;
array2[13647]=30'd611520752;
array2[13648]=30'd611520752;
array2[13649]=30'd611520752;
array2[13650]=30'd611520752;
array2[13651]=30'd611520752;
array2[13652]=30'd611520752;
array2[13653]=30'd606284005;
array2[13654]=30'd611520752;
array2[13655]=30'd611520752;
array2[13656]=30'd611520752;
array2[13657]=30'd611520752;
array2[13658]=30'd606284005;
array2[13659]=30'd611520752;
array2[13660]=30'd606284005;
array2[13661]=30'd611520752;
array2[13662]=30'd606284005;
array2[13663]=30'd611520752;
array2[13664]=30'd611520752;
array2[13665]=30'd611520752;
array2[13666]=30'd611520752;
array2[13667]=30'd611520752;
array2[13668]=30'd611520752;
array2[13669]=30'd611520752;
array2[13670]=30'd611520752;
array2[13671]=30'd619916568;
array2[13672]=30'd401997362;
array2[13673]=30'd865130113;
array2[13674]=30'd851505800;
array2[13675]=30'd851505800;
array2[13676]=30'd858839683;
array2[13677]=30'd858839683;
array2[13678]=30'd851505800;
array2[13679]=30'd851505800;
array2[13680]=30'd858839683;
array2[13681]=30'd865130113;
array2[13682]=30'd858839683;
array2[13683]=30'd858839683;
array2[13684]=30'd858839683;
array2[13685]=30'd858839683;
array2[13686]=30'd858839683;
array2[13687]=30'd851505800;
array2[13688]=30'd858839683;
array2[13689]=30'd858839683;
array2[13690]=30'd858839683;
array2[13691]=30'd851505800;
array2[13692]=30'd858839683;
array2[13693]=30'd858839683;
array2[13694]=30'd865130113;
array2[13695]=30'd858839683;
array2[13696]=30'd858839683;
array2[13697]=30'd858839683;
array2[13698]=30'd865130113;
array2[13699]=30'd858839683;
array2[13700]=30'd858839683;
array2[13701]=30'd799112870;
array2[13702]=30'd718417640;
array2[13703]=30'd732038833;
array2[13704]=30'd851505800;
array2[13705]=30'd851505800;
array2[13706]=30'd858839683;
array2[13707]=30'd819020415;
array2[13708]=30'd770812573;
array2[13709]=30'd606320275;
array2[13710]=30'd347490866;
array2[13711]=30'd240774546;
array2[13712]=30'd227165569;
array2[13713]=30'd227165569;
array2[13714]=30'd234504581;
array2[13715]=30'd230317442;
array2[13716]=30'd231362949;
array2[13717]=30'd231364996;
array2[13718]=30'd231362949;
array2[13719]=30'd231362949;
array2[13720]=30'd229266819;
array2[13721]=30'd229266819;
array2[13722]=30'd231362949;
array2[13723]=30'd231362949;
array2[13724]=30'd234504581;
array2[13725]=30'd231362949;
array2[13726]=30'd231362949;
array2[13727]=30'd231362949;
array2[13728]=30'd559300847;
array2[13729]=30'd595854564;
array2[13730]=30'd595854564;
array2[13731]=30'd606284005;
array2[13732]=30'd586531028;
array2[13733]=30'd586531028;
array2[13734]=30'd586531028;
array2[13735]=30'd586531028;
array2[13736]=30'd586531028;
array2[13737]=30'd586531028;
array2[13738]=30'd586531028;
array2[13739]=30'd586531028;
array2[13740]=30'd586531028;
array2[13741]=30'd586531028;
array2[13742]=30'd585627858;
array2[13743]=30'd586531028;
array2[13744]=30'd595854564;
array2[13745]=30'd595854564;
array2[13746]=30'd595854564;
array2[13747]=30'd595854564;
array2[13748]=30'd595854564;
array2[13749]=30'd595854564;
array2[13750]=30'd595854564;
array2[13751]=30'd595854564;
array2[13752]=30'd595854564;
array2[13753]=30'd595854564;
array2[13754]=30'd611520752;
array2[13755]=30'd586531028;
array2[13756]=30'd586531028;
array2[13757]=30'd586531028;
array2[13758]=30'd586531028;
array2[13759]=30'd586531028;
array2[13760]=30'd586531028;
array2[13761]=30'd586531028;
array2[13762]=30'd586531028;
array2[13763]=30'd586531028;
array2[13764]=30'd586531028;
array2[13765]=30'd585627858;
array2[13766]=30'd586531028;
array2[13767]=30'd582318295;
array2[13768]=30'd401997362;
array2[13769]=30'd865130113;
array2[13770]=30'd851505800;
array2[13771]=30'd851505800;
array2[13772]=30'd858839683;
array2[13773]=30'd858839683;
array2[13774]=30'd858839683;
array2[13775]=30'd851505800;
array2[13776]=30'd858839683;
array2[13777]=30'd858839683;
array2[13778]=30'd858839683;
array2[13779]=30'd858839683;
array2[13780]=30'd858839683;
array2[13781]=30'd851505800;
array2[13782]=30'd858839683;
array2[13783]=30'd851505800;
array2[13784]=30'd858839683;
array2[13785]=30'd851505800;
array2[13786]=30'd858839683;
array2[13787]=30'd851505800;
array2[13788]=30'd858839683;
array2[13789]=30'd858839683;
array2[13790]=30'd858839683;
array2[13791]=30'd858839683;
array2[13792]=30'd858839683;
array2[13793]=30'd858839683;
array2[13794]=30'd851505800;
array2[13795]=30'd858839683;
array2[13796]=30'd851505800;
array2[13797]=30'd865130113;
array2[13798]=30'd865130113;
array2[13799]=30'd851505800;
array2[13800]=30'd858839683;
array2[13801]=30'd851505800;
array2[13802]=30'd770812573;
array2[13803]=30'd713179821;
array2[13804]=30'd560184961;
array2[13805]=30'd260631016;
array2[13806]=30'd240774546;
array2[13807]=30'd262793620;
array2[13808]=30'd238691720;
array2[13809]=30'd238691720;
array2[13810]=30'd227165569;
array2[13811]=30'd231362949;
array2[13812]=30'd231362949;
array2[13813]=30'd231362949;
array2[13814]=30'd231359873;
array2[13815]=30'd231364996;
array2[13816]=30'd231362949;
array2[13817]=30'd229266819;
array2[13818]=30'd231362949;
array2[13819]=30'd231362949;
array2[13820]=30'd231362949;
array2[13821]=30'd231362949;
array2[13822]=30'd231362949;
array2[13823]=30'd229266819;
array2[13824]=30'd498786593;
array2[13825]=30'd543866052;
array2[13826]=30'd561572038;
array2[13827]=30'd561572038;
array2[13828]=30'd537610423;
array2[13829]=30'd530274492;
array2[13830]=30'd530274492;
array2[13831]=30'd537610423;
array2[13832]=30'd530274492;
array2[13833]=30'd530274492;
array2[13834]=30'd514590904;
array2[13835]=30'd530274492;
array2[13836]=30'd530274492;
array2[13837]=30'd514590904;
array2[13838]=30'd524037312;
array2[13839]=30'd537610423;
array2[13840]=30'd543866052;
array2[13841]=30'd543866052;
array2[13842]=30'd543866052;
array2[13843]=30'd543866052;
array2[13844]=30'd543866052;
array2[13845]=30'd543866052;
array2[13846]=30'd543866052;
array2[13847]=30'd543866052;
array2[13848]=30'd543866052;
array2[13849]=30'd543866052;
array2[13850]=30'd561572038;
array2[13851]=30'd543866052;
array2[13852]=30'd530274492;
array2[13853]=30'd530274492;
array2[13854]=30'd530274492;
array2[13855]=30'd530274492;
array2[13856]=30'd530274492;
array2[13857]=30'd537610423;
array2[13858]=30'd530274492;
array2[13859]=30'd530274492;
array2[13860]=30'd530274492;
array2[13861]=30'd514590904;
array2[13862]=30'd530274492;
array2[13863]=30'd561572038;
array2[13864]=30'd401997362;
array2[13865]=30'd865130113;
array2[13866]=30'd858839683;
array2[13867]=30'd858839683;
array2[13868]=30'd858839683;
array2[13869]=30'd851505800;
array2[13870]=30'd858839683;
array2[13871]=30'd851505800;
array2[13872]=30'd858839683;
array2[13873]=30'd851505800;
array2[13874]=30'd865130113;
array2[13875]=30'd858839683;
array2[13876]=30'd858839683;
array2[13877]=30'd851505800;
array2[13878]=30'd851505800;
array2[13879]=30'd851505800;
array2[13880]=30'd858839683;
array2[13881]=30'd858839683;
array2[13882]=30'd858839683;
array2[13883]=30'd858839683;
array2[13884]=30'd858839683;
array2[13885]=30'd858839683;
array2[13886]=30'd858839683;
array2[13887]=30'd851505800;
array2[13888]=30'd851505800;
array2[13889]=30'd770816666;
array2[13890]=30'd713179821;
array2[13891]=30'd770812573;
array2[13892]=30'd799112870;
array2[13893]=30'd770812573;
array2[13894]=30'd770812573;
array2[13895]=30'd770816666;
array2[13896]=30'd770816666;
array2[13897]=30'd732038833;
array2[13898]=30'd601041592;
array2[13899]=30'd347490866;
array2[13900]=30'd281508345;
array2[13901]=30'd248105365;
array2[13902]=30'd240774546;
array2[13903]=30'd227159434;
array2[13904]=30'd234504581;
array2[13905]=30'd234504581;
array2[13906]=30'd234504581;
array2[13907]=30'd231362949;
array2[13908]=30'd230317442;
array2[13909]=30'd231362949;
array2[13910]=30'd231364996;
array2[13911]=30'd231362949;
array2[13912]=30'd228216193;
array2[13913]=30'd231362949;
array2[13914]=30'd231362949;
array2[13915]=30'd234504581;
array2[13916]=30'd231362949;
array2[13917]=30'd234504581;
array2[13918]=30'd231362949;
array2[13919]=30'd231364996;
array2[13920]=30'd496710898;
array2[13921]=30'd518815920;
array2[13922]=30'd518815920;
array2[13923]=30'd518815920;
array2[13924]=30'd518815920;
array2[13925]=30'd518815920;
array2[13926]=30'd518815920;
array2[13927]=30'd518815920;
array2[13928]=30'd518815920;
array2[13929]=30'd518815920;
array2[13930]=30'd518815920;
array2[13931]=30'd518815920;
array2[13932]=30'd518815920;
array2[13933]=30'd518815920;
array2[13934]=30'd518815920;
array2[13935]=30'd521966763;
array2[13936]=30'd521966763;
array2[13937]=30'd518815920;
array2[13938]=30'd518815920;
array2[13939]=30'd518815920;
array2[13940]=30'd518815920;
array2[13941]=30'd518815920;
array2[13942]=30'd518815920;
array2[13943]=30'd518815920;
array2[13944]=30'd518815920;
array2[13945]=30'd518815920;
array2[13946]=30'd518815920;
array2[13947]=30'd518815920;
array2[13948]=30'd518815920;
array2[13949]=30'd518815920;
array2[13950]=30'd518815920;
array2[13951]=30'd521966763;
array2[13952]=30'd521966763;
array2[13953]=30'd518815920;
array2[13954]=30'd521966763;
array2[13955]=30'd518815920;
array2[13956]=30'd518815920;
array2[13957]=30'd521966763;
array2[13958]=30'd518815920;
array2[13959]=30'd514590904;
array2[13960]=30'd401997362;
array2[13961]=30'd828452495;
array2[13962]=30'd851505800;
array2[13963]=30'd858839683;
array2[13964]=30'd858839683;
array2[13965]=30'd858839683;
array2[13966]=30'd858839683;
array2[13967]=30'd851505800;
array2[13968]=30'd851505800;
array2[13969]=30'd858839683;
array2[13970]=30'd865130113;
array2[13971]=30'd858839683;
array2[13972]=30'd858839683;
array2[13973]=30'd858839683;
array2[13974]=30'd858839683;
array2[13975]=30'd858839683;
array2[13976]=30'd858839683;
array2[13977]=30'd865130113;
array2[13978]=30'd858839683;
array2[13979]=30'd858839683;
array2[13980]=30'd858839683;
array2[13981]=30'd858839683;
array2[13982]=30'd858839683;
array2[13983]=30'd858839683;
array2[13984]=30'd851505800;
array2[13985]=30'd770812573;
array2[13986]=30'd606320275;
array2[13987]=30'd560184961;
array2[13988]=30'd678602388;
array2[13989]=30'd711090860;
array2[13990]=30'd678602388;
array2[13991]=30'd672348794;
array2[13992]=30'd606320275;
array2[13993]=30'd401997362;
array2[13994]=30'd281508345;
array2[13995]=30'd228181405;
array2[13996]=30'd265928088;
array2[13997]=30'd262793620;
array2[13998]=30'd238691720;
array2[13999]=30'd262793620;
array2[14000]=30'd234504581;
array2[14001]=30'd231362949;
array2[14002]=30'd229266819;
array2[14003]=30'd231362949;
array2[14004]=30'd229266819;
array2[14005]=30'd231362949;
array2[14006]=30'd229266819;
array2[14007]=30'd229266819;
array2[14008]=30'd229266819;
array2[14009]=30'd229266819;
array2[14010]=30'd230317442;
array2[14011]=30'd229266819;
array2[14012]=30'd229266819;
array2[14013]=30'd229266819;
array2[14014]=30'd231362949;
array2[14015]=30'd227165569;
array2[14016]=30'd496710898;
array2[14017]=30'd518815920;
array2[14018]=30'd524037312;
array2[14019]=30'd518815920;
array2[14020]=30'd515671261;
array2[14021]=30'd515671261;
array2[14022]=30'd520893723;
array2[14023]=30'd515671261;
array2[14024]=30'd515671261;
array2[14025]=30'd515671261;
array2[14026]=30'd515671261;
array2[14027]=30'd515671261;
array2[14028]=30'd515671261;
array2[14029]=30'd515671261;
array2[14030]=30'd510427417;
array2[14031]=30'd515671261;
array2[14032]=30'd521966763;
array2[14033]=30'd518815920;
array2[14034]=30'd515671261;
array2[14035]=30'd518815920;
array2[14036]=30'd518815920;
array2[14037]=30'd518815920;
array2[14038]=30'd518815920;
array2[14039]=30'd518815920;
array2[14040]=30'd521966763;
array2[14041]=30'd515671261;
array2[14042]=30'd518815920;
array2[14043]=30'd521966763;
array2[14044]=30'd515671261;
array2[14045]=30'd515671261;
array2[14046]=30'd515671261;
array2[14047]=30'd515671261;
array2[14048]=30'd515671261;
array2[14049]=30'd515671261;
array2[14050]=30'd515671261;
array2[14051]=30'd515671261;
array2[14052]=30'd515671261;
array2[14053]=30'd510427417;
array2[14054]=30'd515671261;
array2[14055]=30'd518785242;
array2[14056]=30'd381167075;
array2[14057]=30'd727851632;
array2[14058]=30'd851505800;
array2[14059]=30'd865130113;
array2[14060]=30'd858839683;
array2[14061]=30'd858839683;
array2[14062]=30'd858839683;
array2[14063]=30'd865130113;
array2[14064]=30'd865130113;
array2[14065]=30'd865130113;
array2[14066]=30'd858839683;
array2[14067]=30'd858839683;
array2[14068]=30'd858839683;
array2[14069]=30'd858839683;
array2[14070]=30'd858839683;
array2[14071]=30'd858839683;
array2[14072]=30'd858839683;
array2[14073]=30'd828452495;
array2[14074]=30'd828452495;
array2[14075]=30'd828452495;
array2[14076]=30'd805398138;
array2[14077]=30'd805398138;
array2[14078]=30'd828452495;
array2[14079]=30'd828452495;
array2[14080]=30'd819020415;
array2[14081]=30'd819020415;
array2[14082]=30'd672348794;
array2[14083]=30'd483727963;
array2[14084]=30'd481587821;
array2[14085]=30'd485780117;
array2[14086]=30'd407216718;
array2[14087]=30'd178773498;
array2[14088]=30'd190356956;
array2[14089]=30'd254365107;
array2[14090]=30'd262793620;
array2[14091]=30'd262793620;
array2[14092]=30'd262793620;
array2[14093]=30'd262793620;
array2[14094]=30'd238691720;
array2[14095]=30'd238691720;
array2[14096]=30'd234504581;
array2[14097]=30'd234504581;
array2[14098]=30'd231362949;
array2[14099]=30'd231362949;
array2[14100]=30'd231362949;
array2[14101]=30'd231362949;
array2[14102]=30'd229266819;
array2[14103]=30'd230317442;
array2[14104]=30'd231364996;
array2[14105]=30'd231364996;
array2[14106]=30'd229266819;
array2[14107]=30'd228216193;
array2[14108]=30'd229266819;
array2[14109]=30'd229266819;
array2[14110]=30'd231359873;
array2[14111]=30'd234504581;
array2[14112]=30'd387723742;
array2[14113]=30'd475838865;
array2[14114]=30'd475838865;
array2[14115]=30'd475838865;
array2[14116]=30'd477946350;
array2[14117]=30'd477946350;
array2[14118]=30'd477946350;
array2[14119]=30'd477946350;
array2[14120]=30'd477946350;
array2[14121]=30'd477946350;
array2[14122]=30'd473746934;
array2[14123]=30'd477946350;
array2[14124]=30'd473746934;
array2[14125]=30'd477946350;
array2[14126]=30'd477946350;
array2[14127]=30'd477946350;
array2[14128]=30'd475838865;
array2[14129]=30'd475838865;
array2[14130]=30'd475838865;
array2[14131]=30'd475838865;
array2[14132]=30'd475838865;
array2[14133]=30'd475838865;
array2[14134]=30'd475838865;
array2[14135]=30'd475838865;
array2[14136]=30'd477946350;
array2[14137]=30'd475838865;
array2[14138]=30'd475838865;
array2[14139]=30'd477946350;
array2[14140]=30'd477946350;
array2[14141]=30'd477946350;
array2[14142]=30'd477946350;
array2[14143]=30'd477946350;
array2[14144]=30'd477946350;
array2[14145]=30'd477946350;
array2[14146]=30'd477946350;
array2[14147]=30'd477946350;
array2[14148]=30'd477946350;
array2[14149]=30'd473746934;
array2[14150]=30'd473746934;
array2[14151]=30'd475838865;
array2[14152]=30'd387723742;
array2[14153]=30'd450208341;
array2[14154]=30'd828452495;
array2[14155]=30'd858839683;
array2[14156]=30'd858839683;
array2[14157]=30'd851505800;
array2[14158]=30'd858839683;
array2[14159]=30'd858839683;
array2[14160]=30'd858839683;
array2[14161]=30'd851505800;
array2[14162]=30'd858839683;
array2[14163]=30'd858839683;
array2[14164]=30'd851505800;
array2[14165]=30'd858839683;
array2[14166]=30'd828452495;
array2[14167]=30'd828452495;
array2[14168]=30'd799112870;
array2[14169]=30'd770812573;
array2[14170]=30'd732038833;
array2[14171]=30'd732038833;
array2[14172]=30'd601041592;
array2[14173]=30'd678602388;
array2[14174]=30'd732038833;
array2[14175]=30'd770816666;
array2[14176]=30'd819020415;
array2[14177]=30'd819020415;
array2[14178]=30'd768729747;
array2[14179]=30'd566515308;
array2[14180]=30'd481587821;
array2[14181]=30'd539218630;
array2[14182]=30'd434416250;
array2[14183]=30'd179916222;
array2[14184]=30'd238691720;
array2[14185]=30'd238691720;
array2[14186]=30'd238691720;
array2[14187]=30'd238691720;
array2[14188]=30'd238691720;
array2[14189]=30'd238691720;
array2[14190]=30'd238691720;
array2[14191]=30'd234499470;
array2[14192]=30'd227165569;
array2[14193]=30'd234504581;
array2[14194]=30'd234504581;
array2[14195]=30'd231364996;
array2[14196]=30'd231362949;
array2[14197]=30'd230317442;
array2[14198]=30'd229266819;
array2[14199]=30'd231362949;
array2[14200]=30'd231362949;
array2[14201]=30'd231362949;
array2[14202]=30'd231362949;
array2[14203]=30'd231362949;
array2[14204]=30'd231364996;
array2[14205]=30'd231362949;
array2[14206]=30'd231364996;
array2[14207]=30'd231362949;
array2[14208]=30'd439121402;
array2[14209]=30'd482138634;
array2[14210]=30'd482138634;
array2[14211]=30'd475850257;
array2[14212]=30'd482138634;
array2[14213]=30'd475850257;
array2[14214]=30'd475850257;
array2[14215]=30'd482138634;
array2[14216]=30'd482138634;
array2[14217]=30'd475850257;
array2[14218]=30'd482138634;
array2[14219]=30'd482138634;
array2[14220]=30'd475850257;
array2[14221]=30'd475850257;
array2[14222]=30'd482138634;
array2[14223]=30'd482138634;
array2[14224]=30'd482138634;
array2[14225]=30'd475850257;
array2[14226]=30'd482138634;
array2[14227]=30'd475850257;
array2[14228]=30'd475850257;
array2[14229]=30'd482138634;
array2[14230]=30'd482138634;
array2[14231]=30'd475850257;
array2[14232]=30'd480046615;
array2[14233]=30'd480046615;
array2[14234]=30'd475850257;
array2[14235]=30'd482138634;
array2[14236]=30'd482138634;
array2[14237]=30'd475850257;
array2[14238]=30'd480046615;
array2[14239]=30'd480046615;
array2[14240]=30'd482138634;
array2[14241]=30'd482138634;
array2[14242]=30'd475850257;
array2[14243]=30'd480046615;
array2[14244]=30'd480046615;
array2[14245]=30'd480046615;
array2[14246]=30'd482138634;
array2[14247]=30'd490515973;
array2[14248]=30'd439121402;
array2[14249]=30'd425297329;
array2[14250]=30'd606320275;
array2[14251]=30'd828452495;
array2[14252]=30'd851505800;
array2[14253]=30'd858839683;
array2[14254]=30'd858839683;
array2[14255]=30'd858839683;
array2[14256]=30'd858839683;
array2[14257]=30'd858839683;
array2[14258]=30'd851505800;
array2[14259]=30'd851505800;
array2[14260]=30'd828452495;
array2[14261]=30'd770812573;
array2[14262]=30'd732038833;
array2[14263]=30'd732038833;
array2[14264]=30'd732038833;
array2[14265]=30'd604201637;
array2[14266]=30'd407216718;
array2[14267]=30'd407216718;
array2[14268]=30'd347490866;
array2[14269]=30'd347490866;
array2[14270]=30'd606320275;
array2[14271]=30'd711090860;
array2[14272]=30'd768729747;
array2[14273]=30'd819020415;
array2[14274]=30'd819020415;
array2[14275]=30'd678602388;
array2[14276]=30'd506770009;
array2[14277]=30'd539218630;
array2[14278]=30'd434416250;
array2[14279]=30'd179916222;
array2[14280]=30'd238691720;
array2[14281]=30'd228216193;
array2[14282]=30'd231362949;
array2[14283]=30'd228216193;
array2[14284]=30'd229266819;
array2[14285]=30'd231362949;
array2[14286]=30'd228216193;
array2[14287]=30'd230317442;
array2[14288]=30'd231362949;
array2[14289]=30'd229266819;
array2[14290]=30'd229266819;
array2[14291]=30'd229266819;
array2[14292]=30'd231362949;
array2[14293]=30'd231362949;
array2[14294]=30'd231362949;
array2[14295]=30'd230307208;
array2[14296]=30'd229266819;
array2[14297]=30'd230317442;
array2[14298]=30'd231364996;
array2[14299]=30'd229266819;
array2[14300]=30'd229266819;
array2[14301]=30'd228216193;
array2[14302]=30'd229266819;
array2[14303]=30'd229266819;
array2[14304]=30'd387723742;
array2[14305]=30'd457992679;
array2[14306]=30'd473746934;
array2[14307]=30'd490515973;
array2[14308]=30'd457992679;
array2[14309]=30'd439121402;
array2[14310]=30'd439121402;
array2[14311]=30'd439121402;
array2[14312]=30'd439121402;
array2[14313]=30'd439121402;
array2[14314]=30'd439121402;
array2[14315]=30'd457992679;
array2[14316]=30'd439121402;
array2[14317]=30'd439121402;
array2[14318]=30'd387723742;
array2[14319]=30'd457992679;
array2[14320]=30'd473746934;
array2[14321]=30'd473746934;
array2[14322]=30'd473746934;
array2[14323]=30'd490515973;
array2[14324]=30'd473746934;
array2[14325]=30'd473746934;
array2[14326]=30'd473746934;
array2[14327]=30'd473746934;
array2[14328]=30'd457992679;
array2[14329]=30'd473746934;
array2[14330]=30'd475850257;
array2[14331]=30'd457992679;
array2[14332]=30'd457992679;
array2[14333]=30'd457992679;
array2[14334]=30'd439121402;
array2[14335]=30'd439121402;
array2[14336]=30'd439121402;
array2[14337]=30'd439121402;
array2[14338]=30'd439121402;
array2[14339]=30'd457992679;
array2[14340]=30'd439121402;
array2[14341]=30'd387723742;
array2[14342]=30'd439121402;
array2[14343]=30'd509349393;
array2[14344]=30'd457992679;
array2[14345]=30'd528185854;
array2[14346]=30'd425297329;
array2[14347]=30'd678602388;
array2[14348]=30'd770812573;
array2[14349]=30'd851505800;
array2[14350]=30'd858839683;
array2[14351]=30'd865130113;
array2[14352]=30'd858839683;
array2[14353]=30'd851505800;
array2[14354]=30'd851505800;
array2[14355]=30'd828452495;
array2[14356]=30'd764529268;
array2[14357]=30'd606320275;
array2[14358]=30'd713202349;
array2[14359]=30'd678602388;
array2[14360]=30'd450208341;
array2[14361]=30'd319215128;
array2[14362]=30'd193577377;
array2[14363]=30'd212454818;
array2[14364]=30'd212454818;
array2[14365]=30'd186252693;
array2[14366]=30'd319215128;
array2[14367]=30'd606320275;
array2[14368]=30'd713179821;
array2[14369]=30'd819020415;
array2[14370]=30'd819020415;
array2[14371]=30'd805398138;
array2[14372]=30'd483727963;
array2[14373]=30'd539218630;
array2[14374]=30'd281508345;
array2[14375]=30'd232392085;
array2[14376]=30'd232417668;
array2[14377]=30'd229270912;
array2[14378]=30'd231364996;
array2[14379]=30'd231362949;
array2[14380]=30'd231362949;
array2[14381]=30'd231362949;
array2[14382]=30'd228216193;
array2[14383]=30'd229266819;
array2[14384]=30'd231359873;
array2[14385]=30'd231359873;
array2[14386]=30'd231362949;
array2[14387]=30'd234504581;
array2[14388]=30'd231362949;
array2[14389]=30'd231362949;
array2[14390]=30'd230317442;
array2[14391]=30'd229266819;
array2[14392]=30'd229266819;
array2[14393]=30'd229266819;
array2[14394]=30'd230317442;
array2[14395]=30'd230317442;
array2[14396]=30'd230317442;
array2[14397]=30'd228216193;
array2[14398]=30'd231362949;
array2[14399]=30'd234504581;
array2[14400]=30'd307963313;
array2[14401]=30'd340509129;
array2[14402]=30'd340509129;
array2[14403]=30'd340509129;
array2[14404]=30'd307963313;
array2[14405]=30'd302686639;
array2[14406]=30'd302686639;
array2[14407]=30'd302686639;
array2[14408]=30'd302686639;
array2[14409]=30'd302686639;
array2[14410]=30'd302686639;
array2[14411]=30'd302686639;
array2[14412]=30'd302686639;
array2[14413]=30'd265985428;
array2[14414]=30'd232434043;
array2[14415]=30'd302686639;
array2[14416]=30'd340509129;
array2[14417]=30'd362496490;
array2[14418]=30'd340509129;
array2[14419]=30'd340509129;
array2[14420]=30'd340509129;
array2[14421]=30'd340509129;
array2[14422]=30'd340509129;
array2[14423]=30'd340509129;
array2[14424]=30'd340509129;
array2[14425]=30'd340509129;
array2[14426]=30'd340509129;
array2[14427]=30'd307963313;
array2[14428]=30'd302686639;
array2[14429]=30'd302686639;
array2[14430]=30'd302686639;
array2[14431]=30'd302686639;
array2[14432]=30'd302686639;
array2[14433]=30'd302686639;
array2[14434]=30'd302686639;
array2[14435]=30'd302686639;
array2[14436]=30'd265985428;
array2[14437]=30'd235568517;
array2[14438]=30'd302686639;
array2[14439]=30'd362496490;
array2[14440]=30'd307963313;
array2[14441]=30'd362496490;
array2[14442]=30'd302686639;
array2[14443]=30'd518272648;
array2[14444]=30'd711090860;
array2[14445]=30'd770812573;
array2[14446]=30'd828452495;
array2[14447]=30'd851505800;
array2[14448]=30'd851505800;
array2[14449]=30'd819020415;
array2[14450]=30'd819020415;
array2[14451]=30'd819020415;
array2[14452]=30'd805398138;
array2[14453]=30'd646130287;
array2[14454]=30'd383147560;
array2[14455]=30'd281508345;
array2[14456]=30'd207191473;
array2[14457]=30'd213516691;
array2[14458]=30'd227165569;
array2[14459]=30'd234504581;
array2[14460]=30'd231362949;
array2[14461]=30'd228216193;
array2[14462]=30'd220861839;
array2[14463]=30'd347490866;
array2[14464]=30'd604201637;
array2[14465]=30'd768729747;
array2[14466]=30'd819020415;
array2[14467]=30'd819020415;
array2[14468]=30'd483727963;
array2[14469]=30'd450208341;
array2[14470]=30'd179916222;
array2[14471]=30'd231362949;
array2[14472]=30'd229266819;
array2[14473]=30'd229266819;
array2[14474]=30'd229266819;
array2[14475]=30'd228216193;
array2[14476]=30'd228216193;
array2[14477]=30'd230317442;
array2[14478]=30'd230317442;
array2[14479]=30'd229266819;
array2[14480]=30'd234504581;
array2[14481]=30'd229266819;
array2[14482]=30'd234504581;
array2[14483]=30'd231362949;
array2[14484]=30'd231359873;
array2[14485]=30'd231362949;
array2[14486]=30'd230317442;
array2[14487]=30'd229266819;
array2[14488]=30'd230317442;
array2[14489]=30'd228216193;
array2[14490]=30'd228216193;
array2[14491]=30'd230317442;
array2[14492]=30'd229266819;
array2[14493]=30'd229266819;
array2[14494]=30'd231362949;
array2[14495]=30'd231362949;
array2[14496]=30'd193577377;
array2[14497]=30'd228216193;
array2[14498]=30'd227165569;
array2[14499]=30'd227165569;
array2[14500]=30'd228216193;
array2[14501]=30'd228216193;
array2[14502]=30'd232417668;
array2[14503]=30'd234504581;
array2[14504]=30'd231362949;
array2[14505]=30'd229266819;
array2[14506]=30'd229266819;
array2[14507]=30'd227165569;
array2[14508]=30'd231359873;
array2[14509]=30'd230317442;
array2[14510]=30'd231364996;
array2[14511]=30'd231362949;
array2[14512]=30'd234504581;
array2[14513]=30'd228212100;
array2[14514]=30'd228216193;
array2[14515]=30'd229266819;
array2[14516]=30'd231364996;
array2[14517]=30'd228216193;
array2[14518]=30'd228216193;
array2[14519]=30'd231362949;
array2[14520]=30'd229266819;
array2[14521]=30'd231362949;
array2[14522]=30'd228212100;
array2[14523]=30'd227165569;
array2[14524]=30'd231362949;
array2[14525]=30'd231364996;
array2[14526]=30'd234504581;
array2[14527]=30'd234504581;
array2[14528]=30'd234504581;
array2[14529]=30'd227165569;
array2[14530]=30'd231362949;
array2[14531]=30'd228216193;
array2[14532]=30'd234504581;
array2[14533]=30'd262793620;
array2[14534]=30'd240774546;
array2[14535]=30'd257539480;
array2[14536]=30'd262793620;
array2[14537]=30'd265928088;
array2[14538]=30'd257539480;
array2[14539]=30'd260631016;
array2[14540]=30'd407216718;
array2[14541]=30'd711090860;
array2[14542]=30'd799112870;
array2[14543]=30'd819020415;
array2[14544]=30'd819020415;
array2[14545]=30'd819020415;
array2[14546]=30'd819020415;
array2[14547]=30'd819020415;
array2[14548]=30'd805398138;
array2[14549]=30'd645112409;
array2[14550]=30'd207191473;
array2[14551]=30'd227165569;
array2[14552]=30'd230307208;
array2[14553]=30'd231362949;
array2[14554]=30'd229266819;
array2[14555]=30'd229266819;
array2[14556]=30'd228216193;
array2[14557]=30'd230317442;
array2[14558]=30'd229266819;
array2[14559]=30'd228181405;
array2[14560]=30'd383147560;
array2[14561]=30'd711090860;
array2[14562]=30'd805398138;
array2[14563]=30'd805398138;
array2[14564]=30'd444954173;
array2[14565]=30'd179916222;
array2[14566]=30'd227159434;
array2[14567]=30'd234504581;
array2[14568]=30'd229266819;
array2[14569]=30'd229266819;
array2[14570]=30'd231362949;
array2[14571]=30'd231362949;
array2[14572]=30'd231362949;
array2[14573]=30'd231362949;
array2[14574]=30'd231362949;
array2[14575]=30'd229266819;
array2[14576]=30'd231362949;
array2[14577]=30'd231364996;
array2[14578]=30'd234504581;
array2[14579]=30'd231362949;
array2[14580]=30'd231362949;
array2[14581]=30'd231362949;
array2[14582]=30'd230317442;
array2[14583]=30'd229266819;
array2[14584]=30'd229266819;
array2[14585]=30'd231362949;
array2[14586]=30'd231362949;
array2[14587]=30'd231362949;
array2[14588]=30'd231362949;
array2[14589]=30'd234504581;
array2[14590]=30'd231362949;
array2[14591]=30'd228216193;
array2[14592]=30'd193577377;
array2[14593]=30'd227165569;
array2[14594]=30'd227165569;
array2[14595]=30'd231362949;
array2[14596]=30'd234504581;
array2[14597]=30'd231362949;
array2[14598]=30'd231364996;
array2[14599]=30'd228216193;
array2[14600]=30'd231362949;
array2[14601]=30'd231362949;
array2[14602]=30'd231362949;
array2[14603]=30'd231362949;
array2[14604]=30'd228216193;
array2[14605]=30'd229266819;
array2[14606]=30'd231364996;
array2[14607]=30'd231364996;
array2[14608]=30'd231362949;
array2[14609]=30'd231362949;
array2[14610]=30'd231362949;
array2[14611]=30'd231362949;
array2[14612]=30'd231362949;
array2[14613]=30'd234504581;
array2[14614]=30'd228216193;
array2[14615]=30'd234504581;
array2[14616]=30'd229266819;
array2[14617]=30'd229270912;
array2[14618]=30'd228216193;
array2[14619]=30'd234504581;
array2[14620]=30'd228216193;
array2[14621]=30'd234504581;
array2[14622]=30'd227165569;
array2[14623]=30'd234504581;
array2[14624]=30'd231362949;
array2[14625]=30'd231362949;
array2[14626]=30'd229266819;
array2[14627]=30'd231362949;
array2[14628]=30'd240774546;
array2[14629]=30'd265928088;
array2[14630]=30'd262793620;
array2[14631]=30'd262793620;
array2[14632]=30'd265928088;
array2[14633]=30'd262793620;
array2[14634]=30'd262793620;
array2[14635]=30'd265928088;
array2[14636]=30'd260631016;
array2[14637]=30'd401997362;
array2[14638]=30'd672348794;
array2[14639]=30'd768729747;
array2[14640]=30'd805398138;
array2[14641]=30'd819020415;
array2[14642]=30'd819020415;
array2[14643]=30'd805398138;
array2[14644]=30'd713179821;
array2[14645]=30'd565444213;
array2[14646]=30'd207191473;
array2[14647]=30'd231364996;
array2[14648]=30'd231364996;
array2[14649]=30'd231364996;
array2[14650]=30'd229266819;
array2[14651]=30'd231362949;
array2[14652]=30'd228216193;
array2[14653]=30'd229266819;
array2[14654]=30'd229266819;
array2[14655]=30'd220861839;
array2[14656]=30'd281508345;
array2[14657]=30'd560184961;
array2[14658]=30'd711090860;
array2[14659]=30'd631447172;
array2[14660]=30'd260631016;
array2[14661]=30'd227165569;
array2[14662]=30'd231362949;
array2[14663]=30'd230317442;
array2[14664]=30'd231364996;
array2[14665]=30'd231362949;
array2[14666]=30'd231362949;
array2[14667]=30'd228216193;
array2[14668]=30'd228216193;
array2[14669]=30'd229266819;
array2[14670]=30'd231362949;
array2[14671]=30'd231359873;
array2[14672]=30'd231362949;
array2[14673]=30'd234504581;
array2[14674]=30'd231362949;
array2[14675]=30'd231364996;
array2[14676]=30'd231364996;
array2[14677]=30'd229266819;
array2[14678]=30'd229266819;
array2[14679]=30'd229266819;
array2[14680]=30'd230317442;
array2[14681]=30'd230317442;
array2[14682]=30'd230317442;
array2[14683]=30'd228216193;
array2[14684]=30'd228216193;
array2[14685]=30'd234504581;
array2[14686]=30'd231362949;
array2[14687]=30'd231362949;
array2[14688]=30'd212454818;
array2[14689]=30'd234504581;
array2[14690]=30'd228212100;
array2[14691]=30'd230317442;
array2[14692]=30'd230317442;
array2[14693]=30'd230317442;
array2[14694]=30'd231362949;
array2[14695]=30'd230317442;
array2[14696]=30'd231362949;
array2[14697]=30'd231362949;
array2[14698]=30'd231362949;
array2[14699]=30'd231362949;
array2[14700]=30'd231362949;
array2[14701]=30'd229266819;
array2[14702]=30'd231362949;
array2[14703]=30'd234504581;
array2[14704]=30'd231364996;
array2[14705]=30'd229266819;
array2[14706]=30'd229266819;
array2[14707]=30'd231362949;
array2[14708]=30'd231362949;
array2[14709]=30'd231362949;
array2[14710]=30'd231362949;
array2[14711]=30'd231362949;
array2[14712]=30'd231362949;
array2[14713]=30'd231364996;
array2[14714]=30'd229270912;
array2[14715]=30'd234504581;
array2[14716]=30'd231362949;
array2[14717]=30'd234504581;
array2[14718]=30'd231362949;
array2[14719]=30'd230317442;
array2[14720]=30'd228216193;
array2[14721]=30'd228216193;
array2[14722]=30'd231359873;
array2[14723]=30'd232392085;
array2[14724]=30'd265928088;
array2[14725]=30'd265928088;
array2[14726]=30'd238691720;
array2[14727]=30'd234504581;
array2[14728]=30'd234504581;
array2[14729]=30'd234504581;
array2[14730]=30'd238691720;
array2[14731]=30'd234504581;
array2[14732]=30'd227159434;
array2[14733]=30'd190356956;
array2[14734]=30'd401997362;
array2[14735]=30'd672348794;
array2[14736]=30'd768729747;
array2[14737]=30'd819020415;
array2[14738]=30'd805398138;
array2[14739]=30'd768729747;
array2[14740]=30'd606320275;
array2[14741]=30'd383147560;
array2[14742]=30'd228181405;
array2[14743]=30'd231362949;
array2[14744]=30'd231364996;
array2[14745]=30'd229266819;
array2[14746]=30'd229266819;
array2[14747]=30'd231362949;
array2[14748]=30'd231362949;
array2[14749]=30'd231362949;
array2[14750]=30'd231362949;
array2[14751]=30'd231359873;
array2[14752]=30'd228181405;
array2[14753]=30'd338018898;
array2[14754]=30'd565444213;
array2[14755]=30'd347490866;
array2[14756]=30'd232392085;
array2[14757]=30'd231362949;
array2[14758]=30'd231362949;
array2[14759]=30'd229266819;
array2[14760]=30'd231364996;
array2[14761]=30'd228216193;
array2[14762]=30'd228216193;
array2[14763]=30'd229266819;
array2[14764]=30'd230317442;
array2[14765]=30'd229266819;
array2[14766]=30'd234504581;
array2[14767]=30'd231359873;
array2[14768]=30'd231362949;
array2[14769]=30'd231362949;
array2[14770]=30'd229266819;
array2[14771]=30'd231362949;
array2[14772]=30'd231362949;
array2[14773]=30'd231362949;
array2[14774]=30'd229266819;
array2[14775]=30'd229266819;
array2[14776]=30'd231362949;
array2[14777]=30'd231364996;
array2[14778]=30'd229270912;
array2[14779]=30'd231359873;
array2[14780]=30'd234504581;
array2[14781]=30'd231362949;
array2[14782]=30'd231362949;
array2[14783]=30'd229270912;
array2[14784]=30'd212454818;
array2[14785]=30'd234504581;
array2[14786]=30'd228212100;
array2[14787]=30'd230317442;
array2[14788]=30'd230317442;
array2[14789]=30'd230317442;
array2[14790]=30'd231362949;
array2[14791]=30'd230317442;
array2[14792]=30'd231362949;
array2[14793]=30'd231362949;
array2[14794]=30'd231362949;
array2[14795]=30'd231362949;
array2[14796]=30'd231362949;
array2[14797]=30'd229266819;
array2[14798]=30'd231362949;
array2[14799]=30'd234504581;
array2[14800]=30'd231359873;
array2[14801]=30'd231364996;
array2[14802]=30'd229266819;
array2[14803]=30'd229266819;
array2[14804]=30'd231362949;
array2[14805]=30'd228216193;
array2[14806]=30'd231362949;
array2[14807]=30'd231362949;
array2[14808]=30'd231362949;
array2[14809]=30'd231362949;
array2[14810]=30'd231364996;
array2[14811]=30'd231364996;
array2[14812]=30'd234504581;
array2[14813]=30'd231362949;
array2[14814]=30'd234504581;
array2[14815]=30'd231364996;
array2[14816]=30'd230317442;
array2[14817]=30'd229266819;
array2[14818]=30'd228216193;
array2[14819]=30'd238691720;
array2[14820]=30'd262793620;
array2[14821]=30'd227165569;
array2[14822]=30'd236604812;
array2[14823]=30'd231364996;
array2[14824]=30'd231362949;
array2[14825]=30'd229266819;
array2[14826]=30'd231362949;
array2[14827]=30'd231362949;
array2[14828]=30'd230307208;
array2[14829]=30'd190356956;
array2[14830]=30'd338018898;
array2[14831]=30'd506770009;
array2[14832]=30'd678602388;
array2[14833]=30'd805398138;
array2[14834]=30'd711090860;
array2[14835]=30'd481587821;
array2[14836]=30'd347490866;
array2[14837]=30'd212454818;
array2[14838]=30'd227165569;
array2[14839]=30'd231362949;
array2[14840]=30'd231362949;
array2[14841]=30'd229266819;
array2[14842]=30'd231362949;
array2[14843]=30'd234504581;
array2[14844]=30'd229266819;
array2[14845]=30'd229266819;
array2[14846]=30'd231362949;
array2[14847]=30'd231362949;
array2[14848]=30'd265928088;
array2[14849]=30'd260631016;
array2[14850]=30'd260631016;
array2[14851]=30'd260631016;
array2[14852]=30'd221916546;
array2[14853]=30'd229266819;
array2[14854]=30'd231362949;
array2[14855]=30'd230317442;
array2[14856]=30'd230317442;
array2[14857]=30'd231362949;
array2[14858]=30'd231362949;
array2[14859]=30'd231362949;
array2[14860]=30'd229266819;
array2[14861]=30'd231362949;
array2[14862]=30'd231362949;
array2[14863]=30'd231362949;
array2[14864]=30'd231362949;
array2[14865]=30'd231362949;
array2[14866]=30'd230317442;
array2[14867]=30'd231362949;
array2[14868]=30'd230317442;
array2[14869]=30'd229266819;
array2[14870]=30'd229266819;
array2[14871]=30'd229266819;
array2[14872]=30'd231364996;
array2[14873]=30'd229266819;
array2[14874]=30'd231362949;
array2[14875]=30'd234504581;
array2[14876]=30'd231362949;
array2[14877]=30'd234504581;
array2[14878]=30'd230317442;
array2[14879]=30'd229266819;
array2[14880]=30'd193577377;
array2[14881]=30'd227165569;
array2[14882]=30'd228212100;
array2[14883]=30'd231362949;
array2[14884]=30'd231362949;
array2[14885]=30'd231362949;
array2[14886]=30'd231364996;
array2[14887]=30'd229266819;
array2[14888]=30'd231364996;
array2[14889]=30'd231362949;
array2[14890]=30'd231362949;
array2[14891]=30'd231362949;
array2[14892]=30'd231362949;
array2[14893]=30'd229266819;
array2[14894]=30'd231362949;
array2[14895]=30'd234504581;
array2[14896]=30'd231362949;
array2[14897]=30'd231364996;
array2[14898]=30'd231364996;
array2[14899]=30'd231362949;
array2[14900]=30'd231362949;
array2[14901]=30'd228216193;
array2[14902]=30'd229266819;
array2[14903]=30'd229266819;
array2[14904]=30'd231362949;
array2[14905]=30'd231362949;
array2[14906]=30'd231362949;
array2[14907]=30'd231362949;
array2[14908]=30'd231362949;
array2[14909]=30'd231362949;
array2[14910]=30'd231364996;
array2[14911]=30'd231362949;
array2[14912]=30'd229266819;
array2[14913]=30'd229266819;
array2[14914]=30'd230317442;
array2[14915]=30'd231362949;
array2[14916]=30'd238691720;
array2[14917]=30'd231362949;
array2[14918]=30'd231362949;
array2[14919]=30'd231362949;
array2[14920]=30'd231362949;
array2[14921]=30'd231362949;
array2[14922]=30'd231362949;
array2[14923]=30'd230317442;
array2[14924]=30'd231362949;
array2[14925]=30'd228181405;
array2[14926]=30'd319215128;
array2[14927]=30'd450208341;
array2[14928]=30'd560184961;
array2[14929]=30'd768729747;
array2[14930]=30'd764529268;
array2[14931]=30'd450208341;
array2[14932]=30'd383147560;
array2[14933]=30'd238691720;
array2[14934]=30'd228216193;
array2[14935]=30'd229270912;
array2[14936]=30'd228216193;
array2[14937]=30'd231359873;
array2[14938]=30'd231364996;
array2[14939]=30'd229266819;
array2[14940]=30'd229266819;
array2[14941]=30'd231362949;
array2[14942]=30'd231359873;
array2[14943]=30'd231362949;
array2[14944]=30'd231362949;
array2[14945]=30'd231362949;
array2[14946]=30'd229266819;
array2[14947]=30'd229270912;
array2[14948]=30'd231364996;
array2[14949]=30'd234504581;
array2[14950]=30'd231362949;
array2[14951]=30'd231362949;
array2[14952]=30'd231364996;
array2[14953]=30'd230317442;
array2[14954]=30'd229266819;
array2[14955]=30'd228216193;
array2[14956]=30'd231362949;
array2[14957]=30'd231362949;
array2[14958]=30'd231362949;
array2[14959]=30'd231362949;
array2[14960]=30'd234504581;
array2[14961]=30'd231362949;
array2[14962]=30'd227165569;
array2[14963]=30'd227165569;
array2[14964]=30'd231364996;
array2[14965]=30'd230317442;
array2[14966]=30'd231362949;
array2[14967]=30'd231362949;
array2[14968]=30'd231364996;
array2[14969]=30'd231362949;
array2[14970]=30'd231362949;
array2[14971]=30'd231362949;
array2[14972]=30'd234504581;
array2[14973]=30'd229266819;
array2[14974]=30'd231362949;
array2[14975]=30'd231364996;
array2[14976]=30'd193577377;
array2[14977]=30'd227165569;
array2[14978]=30'd228212100;
array2[14979]=30'd231362949;
array2[14980]=30'd231362949;
array2[14981]=30'd231362949;
array2[14982]=30'd231364996;
array2[14983]=30'd229266819;
array2[14984]=30'd231362949;
array2[14985]=30'd231362949;
array2[14986]=30'd231362949;
array2[14987]=30'd231362949;
array2[14988]=30'd228216193;
array2[14989]=30'd229266819;
array2[14990]=30'd231362949;
array2[14991]=30'd234504581;
array2[14992]=30'd231362949;
array2[14993]=30'd231362949;
array2[14994]=30'd230317442;
array2[14995]=30'd231362949;
array2[14996]=30'd231362949;
array2[14997]=30'd231362949;
array2[14998]=30'd228216193;
array2[14999]=30'd228216193;
array2[15000]=30'd229266819;
array2[15001]=30'd231362949;
array2[15002]=30'd231364996;
array2[15003]=30'd231359873;
array2[15004]=30'd231364996;
array2[15005]=30'd231362949;
array2[15006]=30'd230317442;
array2[15007]=30'd231362949;
array2[15008]=30'd229266819;
array2[15009]=30'd228216193;
array2[15010]=30'd229266819;
array2[15011]=30'd231364996;
array2[15012]=30'd231364996;
array2[15013]=30'd230317442;
array2[15014]=30'd231362949;
array2[15015]=30'd234504581;
array2[15016]=30'd230317442;
array2[15017]=30'd231362949;
array2[15018]=30'd229266819;
array2[15019]=30'd229266819;
array2[15020]=30'd231364996;
array2[15021]=30'd228216193;
array2[15022]=30'd228181405;
array2[15023]=30'd249001484;
array2[15024]=30'd249001484;
array2[15025]=30'd566515308;
array2[15026]=30'd678602388;
array2[15027]=30'd672348794;
array2[15028]=30'd560184961;
array2[15029]=30'd381167075;
array2[15030]=30'd234504581;
array2[15031]=30'd232417668;
array2[15032]=30'd231364996;
array2[15033]=30'd231359873;
array2[15034]=30'd231364996;
array2[15035]=30'd229266819;
array2[15036]=30'd229266819;
array2[15037]=30'd231362949;
array2[15038]=30'd231362949;
array2[15039]=30'd231362949;
array2[15040]=30'd231362949;
array2[15041]=30'd231362949;
array2[15042]=30'd231362949;
array2[15043]=30'd231364996;
array2[15044]=30'd231364996;
array2[15045]=30'd234504581;
array2[15046]=30'd231362949;
array2[15047]=30'd231362949;
array2[15048]=30'd231362949;
array2[15049]=30'd230317442;
array2[15050]=30'd228216193;
array2[15051]=30'd228216193;
array2[15052]=30'd231362949;
array2[15053]=30'd231362949;
array2[15054]=30'd231362949;
array2[15055]=30'd231362949;
array2[15056]=30'd234504581;
array2[15057]=30'd228216193;
array2[15058]=30'd234504581;
array2[15059]=30'd227165569;
array2[15060]=30'd231362949;
array2[15061]=30'd230317442;
array2[15062]=30'd230317442;
array2[15063]=30'd231364996;
array2[15064]=30'd231362949;
array2[15065]=30'd228216193;
array2[15066]=30'd228216193;
array2[15067]=30'd229266819;
array2[15068]=30'd229266819;
array2[15069]=30'd231362949;
array2[15070]=30'd231362949;
array2[15071]=30'd234504581;
array2[15072]=30'd193577377;
array2[15073]=30'd227165569;
array2[15074]=30'd228212100;
array2[15075]=30'd231362949;
array2[15076]=30'd231362949;
array2[15077]=30'd231362949;
array2[15078]=30'd231364996;
array2[15079]=30'd229266819;
array2[15080]=30'd231362949;
array2[15081]=30'd231362949;
array2[15082]=30'd229266819;
array2[15083]=30'd229266819;
array2[15084]=30'd228216193;
array2[15085]=30'd230317442;
array2[15086]=30'd231362949;
array2[15087]=30'd231362949;
array2[15088]=30'd231362949;
array2[15089]=30'd229266819;
array2[15090]=30'd231359873;
array2[15091]=30'd231364996;
array2[15092]=30'd231362949;
array2[15093]=30'd229266819;
array2[15094]=30'd234504581;
array2[15095]=30'd231362949;
array2[15096]=30'd231362949;
array2[15097]=30'd229266819;
array2[15098]=30'd231362949;
array2[15099]=30'd231362949;
array2[15100]=30'd231364996;
array2[15101]=30'd231364996;
array2[15102]=30'd231359873;
array2[15103]=30'd231362949;
array2[15104]=30'd231362949;
array2[15105]=30'd231364996;
array2[15106]=30'd230317442;
array2[15107]=30'd231362949;
array2[15108]=30'd228216193;
array2[15109]=30'd231362949;
array2[15110]=30'd231362949;
array2[15111]=30'd229266819;
array2[15112]=30'd231362949;
array2[15113]=30'd231362949;
array2[15114]=30'd231362949;
array2[15115]=30'd234504581;
array2[15116]=30'd228216193;
array2[15117]=30'd231364996;
array2[15118]=30'd228216193;
array2[15119]=30'd220861839;
array2[15120]=30'd195647926;
array2[15121]=30'd249001484;
array2[15122]=30'd319215128;
array2[15123]=30'd319215128;
array2[15124]=30'd281508345;
array2[15125]=30'd190356956;
array2[15126]=30'd212454818;
array2[15127]=30'd227165569;
array2[15128]=30'd228216193;
array2[15129]=30'd231362949;
array2[15130]=30'd231362949;
array2[15131]=30'd228216193;
array2[15132]=30'd229270912;
array2[15133]=30'd231362949;
array2[15134]=30'd231362949;
array2[15135]=30'd231359873;
array2[15136]=30'd230317442;
array2[15137]=30'd231362949;
array2[15138]=30'd229266819;
array2[15139]=30'd231362949;
array2[15140]=30'd231359873;
array2[15141]=30'd231362949;
array2[15142]=30'd231364996;
array2[15143]=30'd229266819;
array2[15144]=30'd229266819;
array2[15145]=30'd231364996;
array2[15146]=30'd231362949;
array2[15147]=30'd231362949;
array2[15148]=30'd229266819;
array2[15149]=30'd234504581;
array2[15150]=30'd231362949;
array2[15151]=30'd229266819;
array2[15152]=30'd228216193;
array2[15153]=30'd228216193;
array2[15154]=30'd228216193;
array2[15155]=30'd231364996;
array2[15156]=30'd231362949;
array2[15157]=30'd231362949;
array2[15158]=30'd231362949;
array2[15159]=30'd229266819;
array2[15160]=30'd228216193;
array2[15161]=30'd227165569;
array2[15162]=30'd231364996;
array2[15163]=30'd229266819;
array2[15164]=30'd228216193;
array2[15165]=30'd231362949;
array2[15166]=30'd230317442;
array2[15167]=30'd229266819;
array2[15168]=30'd193577377;
array2[15169]=30'd227165569;
array2[15170]=30'd227165569;
array2[15171]=30'd272255371;
array2[15172]=30'd236604812;
array2[15173]=30'd231362949;
array2[15174]=30'd231362949;
array2[15175]=30'd229266819;
array2[15176]=30'd229266819;
array2[15177]=30'd231362949;
array2[15178]=30'd231362949;
array2[15179]=30'd231362949;
array2[15180]=30'd231362949;
array2[15181]=30'd234504581;
array2[15182]=30'd301610387;
array2[15183]=30'd256519562;
array2[15184]=30'd231362949;
array2[15185]=30'd231362949;
array2[15186]=30'd231364996;
array2[15187]=30'd230317442;
array2[15188]=30'd229266819;
array2[15189]=30'd231362949;
array2[15190]=30'd231362949;
array2[15191]=30'd228216193;
array2[15192]=30'd229266819;
array2[15193]=30'd229266819;
array2[15194]=30'd256519562;
array2[15195]=30'd256519562;
array2[15196]=30'd231362949;
array2[15197]=30'd231362949;
array2[15198]=30'd230317442;
array2[15199]=30'd230317442;
array2[15200]=30'd231364996;
array2[15201]=30'd229266819;
array2[15202]=30'd228216193;
array2[15203]=30'd231362949;
array2[15204]=30'd229266819;
array2[15205]=30'd338288022;
array2[15206]=30'd272255371;
array2[15207]=30'd230307208;
array2[15208]=30'd231359873;
array2[15209]=30'd229266819;
array2[15210]=30'd231362949;
array2[15211]=30'd229266819;
array2[15212]=30'd229266819;
array2[15213]=30'd229266819;
array2[15214]=30'd231364996;
array2[15215]=30'd230317442;
array2[15216]=30'd230307208;
array2[15217]=30'd227159434;
array2[15218]=30'd227159434;
array2[15219]=30'd227159434;
array2[15220]=30'd227159434;
array2[15221]=30'd227159434;
array2[15222]=30'd227165569;
array2[15223]=30'd229266819;
array2[15224]=30'd229266819;
array2[15225]=30'd229266819;
array2[15226]=30'd231362949;
array2[15227]=30'd231362949;
array2[15228]=30'd231362949;
array2[15229]=30'd230317442;
array2[15230]=30'd230317442;
array2[15231]=30'd229266819;
array2[15232]=30'd229266819;
array2[15233]=30'd231362949;
array2[15234]=30'd231362949;
array2[15235]=30'd229266819;
array2[15236]=30'd229266819;
array2[15237]=30'd228216193;
array2[15238]=30'd231364996;
array2[15239]=30'd229266819;
array2[15240]=30'd229266819;
array2[15241]=30'd229266819;
array2[15242]=30'd229266819;
array2[15243]=30'd231362949;
array2[15244]=30'd229266819;
array2[15245]=30'd230317442;
array2[15246]=30'd231362949;
array2[15247]=30'd229266819;
array2[15248]=30'd231362949;
array2[15249]=30'd229266819;
array2[15250]=30'd231362949;
array2[15251]=30'd231362949;
array2[15252]=30'd231362949;
array2[15253]=30'd230317442;
array2[15254]=30'd230317442;
array2[15255]=30'd229266819;
array2[15256]=30'd231362949;
array2[15257]=30'd231362949;
array2[15258]=30'd234504581;
array2[15259]=30'd229266819;
array2[15260]=30'd229266819;
array2[15261]=30'd231362949;
array2[15262]=30'd229266819;
array2[15263]=30'd231362949;
array2[15264]=30'd193577377;
array2[15265]=30'd230307208;
array2[15266]=30'd272255371;
array2[15267]=30'd472496545;
array2[15268]=30'd272255371;
array2[15269]=30'd229266819;
array2[15270]=30'd231364996;
array2[15271]=30'd229266819;
array2[15272]=30'd231364996;
array2[15273]=30'd231362949;
array2[15274]=30'd231362949;
array2[15275]=30'd256519562;
array2[15276]=30'd236604812;
array2[15277]=30'd272255371;
array2[15278]=30'd710509991;
array2[15279]=30'd425297329;
array2[15280]=30'd234499470;
array2[15281]=30'd256519562;
array2[15282]=30'd234504581;
array2[15283]=30'd228216193;
array2[15284]=30'd231359873;
array2[15285]=30'd231362949;
array2[15286]=30'd231362949;
array2[15287]=30'd231362949;
array2[15288]=30'd229266819;
array2[15289]=30'd231362949;
array2[15290]=30'd472496545;
array2[15291]=30'd338288022;
array2[15292]=30'd230317442;
array2[15293]=30'd231364996;
array2[15294]=30'd229266819;
array2[15295]=30'd231362949;
array2[15296]=30'd231362949;
array2[15297]=30'd231362949;
array2[15298]=30'd238691720;
array2[15299]=30'd238691720;
array2[15300]=30'd256519562;
array2[15301]=30'd655981997;
array2[15302]=30'd472496545;
array2[15303]=30'd221916546;
array2[15304]=30'd272255371;
array2[15305]=30'd230307208;
array2[15306]=30'd231362949;
array2[15307]=30'd231364996;
array2[15308]=30'd230317442;
array2[15309]=30'd228216193;
array2[15310]=30'd228216193;
array2[15311]=30'd231362949;
array2[15312]=30'd230317442;
array2[15313]=30'd229266819;
array2[15314]=30'd234504581;
array2[15315]=30'd234504581;
array2[15316]=30'd231359873;
array2[15317]=30'd230317442;
array2[15318]=30'd229266819;
array2[15319]=30'd229266819;
array2[15320]=30'd231362949;
array2[15321]=30'd231362949;
array2[15322]=30'd231362949;
array2[15323]=30'd231362949;
array2[15324]=30'd231362949;
array2[15325]=30'd227165569;
array2[15326]=30'd231364996;
array2[15327]=30'd231362949;
array2[15328]=30'd234504581;
array2[15329]=30'd231362949;
array2[15330]=30'd231362949;
array2[15331]=30'd231362949;
array2[15332]=30'd231362949;
array2[15333]=30'd229266819;
array2[15334]=30'd229266819;
array2[15335]=30'd231362949;
array2[15336]=30'd231362949;
array2[15337]=30'd229266819;
array2[15338]=30'd231362949;
array2[15339]=30'd231362949;
array2[15340]=30'd229266819;
array2[15341]=30'd230307208;
array2[15342]=30'd227165569;
array2[15343]=30'd231364996;
array2[15344]=30'd230317442;
array2[15345]=30'd231362949;
array2[15346]=30'd231364996;
array2[15347]=30'd231364996;
array2[15348]=30'd231362949;
array2[15349]=30'd231362949;
array2[15350]=30'd229266819;
array2[15351]=30'd231362949;
array2[15352]=30'd231362949;
array2[15353]=30'd231362949;
array2[15354]=30'd234504581;
array2[15355]=30'd231362949;
array2[15356]=30'd231362949;
array2[15357]=30'd231362949;
array2[15358]=30'd231362949;
array2[15359]=30'd229266819;
array2[15360]=30'd193577377;
array2[15361]=30'd227165569;
array2[15362]=30'd272255371;
array2[15363]=30'd472496545;
array2[15364]=30'd272255371;
array2[15365]=30'd228216193;
array2[15366]=30'd231359873;
array2[15367]=30'd231362949;
array2[15368]=30'd230317442;
array2[15369]=30'd231362949;
array2[15370]=30'd231362949;
array2[15371]=30'd664345022;
array2[15372]=30'd425297329;
array2[15373]=30'd238691720;
array2[15374]=30'd272255371;
array2[15375]=30'd256519562;
array2[15376]=30'd377085336;
array2[15377]=30'd664345022;
array2[15378]=30'd256519562;
array2[15379]=30'd231364996;
array2[15380]=30'd231362949;
array2[15381]=30'd230317442;
array2[15382]=30'd231362949;
array2[15383]=30'd229266819;
array2[15384]=30'd231362949;
array2[15385]=30'd231362949;
array2[15386]=30'd428475791;
array2[15387]=30'd338288022;
array2[15388]=30'd230307208;
array2[15389]=30'd229266819;
array2[15390]=30'd231364996;
array2[15391]=30'd231362949;
array2[15392]=30'd229266819;
array2[15393]=30'd227165569;
array2[15394]=30'd532258209;
array2[15395]=30'd553231776;
array2[15396]=30'd227165569;
array2[15397]=30'd272255371;
array2[15398]=30'd256519562;
array2[15399]=30'd256519562;
array2[15400]=30'd655981997;
array2[15401]=30'd281654691;
array2[15402]=30'd234504581;
array2[15403]=30'd229266819;
array2[15404]=30'd231362949;
array2[15405]=30'd231362949;
array2[15406]=30'd230317442;
array2[15407]=30'd228216193;
array2[15408]=30'd231362949;
array2[15409]=30'd231362949;
array2[15410]=30'd231359873;
array2[15411]=30'd231362949;
array2[15412]=30'd231359873;
array2[15413]=30'd230317442;
array2[15414]=30'd231364996;
array2[15415]=30'd230317442;
array2[15416]=30'd234504581;
array2[15417]=30'd231362949;
array2[15418]=30'd231362949;
array2[15419]=30'd231362949;
array2[15420]=30'd230317442;
array2[15421]=30'd228216193;
array2[15422]=30'd230317442;
array2[15423]=30'd231362949;
array2[15424]=30'd231362949;
array2[15425]=30'd231362949;
array2[15426]=30'd234504581;
array2[15427]=30'd231362949;
array2[15428]=30'd231362949;
array2[15429]=30'd228216193;
array2[15430]=30'd227165569;
array2[15431]=30'd231362949;
array2[15432]=30'd231362949;
array2[15433]=30'd228216193;
array2[15434]=30'd231362949;
array2[15435]=30'd234504581;
array2[15436]=30'd231362949;
array2[15437]=30'd228216193;
array2[15438]=30'd227165569;
array2[15439]=30'd231364996;
array2[15440]=30'd231362949;
array2[15441]=30'd234504581;
array2[15442]=30'd231362949;
array2[15443]=30'd231362949;
array2[15444]=30'd231362949;
array2[15445]=30'd231362949;
array2[15446]=30'd231364996;
array2[15447]=30'd234504581;
array2[15448]=30'd231362949;
array2[15449]=30'd231362949;
array2[15450]=30'd231364996;
array2[15451]=30'd231364996;
array2[15452]=30'd229266819;
array2[15453]=30'd229266819;
array2[15454]=30'd231362949;
array2[15455]=30'd231362949;
array2[15456]=30'd212454818;
array2[15457]=30'd238691720;
array2[15458]=30'd227165569;
array2[15459]=30'd256519562;
array2[15460]=30'd234504581;
array2[15461]=30'd227165569;
array2[15462]=30'd234504581;
array2[15463]=30'd234504581;
array2[15464]=30'd234504581;
array2[15465]=30'd231364996;
array2[15466]=30'd256519562;
array2[15467]=30'd262793620;
array2[15468]=30'd236604812;
array2[15469]=30'd234504581;
array2[15470]=30'd231364996;
array2[15471]=30'd231364996;
array2[15472]=30'd236604812;
array2[15473]=30'd256519562;
array2[15474]=30'd256519562;
array2[15475]=30'd229270912;
array2[15476]=30'd231364996;
array2[15477]=30'd231362949;
array2[15478]=30'd234504581;
array2[15479]=30'd229266819;
array2[15480]=30'd231362949;
array2[15481]=30'd231362949;
array2[15482]=30'd256519562;
array2[15483]=30'd232417668;
array2[15484]=30'd234504581;
array2[15485]=30'd231359873;
array2[15486]=30'd234504581;
array2[15487]=30'd229266819;
array2[15488]=30'd234504581;
array2[15489]=30'd256519562;
array2[15490]=30'd256519562;
array2[15491]=30'd256519562;
array2[15492]=30'd231362949;
array2[15493]=30'd229266819;
array2[15494]=30'd231364996;
array2[15495]=30'd228216193;
array2[15496]=30'd256519562;
array2[15497]=30'd234504581;
array2[15498]=30'd256519562;
array2[15499]=30'd228216193;
array2[15500]=30'd234504581;
array2[15501]=30'd229266819;
array2[15502]=30'd229266819;
array2[15503]=30'd231362949;
array2[15504]=30'd228216193;
array2[15505]=30'd231362949;
array2[15506]=30'd231362949;
array2[15507]=30'd229266819;
array2[15508]=30'd229266819;
array2[15509]=30'd231362949;
array2[15510]=30'd231359873;
array2[15511]=30'd229266819;
array2[15512]=30'd231362949;
array2[15513]=30'd231362949;
array2[15514]=30'd229266819;
array2[15515]=30'd230317442;
array2[15516]=30'd229266819;
array2[15517]=30'd231362949;
array2[15518]=30'd230317442;
array2[15519]=30'd234504581;
array2[15520]=30'd228216193;
array2[15521]=30'd229266819;
array2[15522]=30'd230317442;
array2[15523]=30'd231364996;
array2[15524]=30'd229266819;
array2[15525]=30'd231359873;
array2[15526]=30'd231362949;
array2[15527]=30'd230317442;
array2[15528]=30'd231364996;
array2[15529]=30'd231362949;
array2[15530]=30'd231362949;
array2[15531]=30'd228216193;
array2[15532]=30'd231362949;
array2[15533]=30'd229266819;
array2[15534]=30'd230317442;
array2[15535]=30'd229266819;
array2[15536]=30'd231362949;
array2[15537]=30'd231364996;
array2[15538]=30'd231362949;
array2[15539]=30'd231362949;
array2[15540]=30'd231362949;
array2[15541]=30'd229266819;
array2[15542]=30'd229266819;
array2[15543]=30'd231362949;
array2[15544]=30'd231362949;
array2[15545]=30'd231364996;
array2[15546]=30'd231364996;
array2[15547]=30'd231362949;
array2[15548]=30'd228216193;
array2[15549]=30'd231362949;
array2[15550]=30'd231362949;
array2[15551]=30'd229266819;
array2[15552]=30'd212454818;
array2[15553]=30'd234504581;
array2[15554]=30'd227165569;
array2[15555]=30'd231362949;
array2[15556]=30'd234504581;
array2[15557]=30'd229266819;
array2[15558]=30'd231362949;
array2[15559]=30'd231362949;
array2[15560]=30'd231364996;
array2[15561]=30'd229266819;
array2[15562]=30'd234504581;
array2[15563]=30'd234504581;
array2[15564]=30'd231362949;
array2[15565]=30'd231364996;
array2[15566]=30'd230317442;
array2[15567]=30'd229266819;
array2[15568]=30'd229266819;
array2[15569]=30'd231362949;
array2[15570]=30'd234504581;
array2[15571]=30'd227165569;
array2[15572]=30'd234504581;
array2[15573]=30'd234504581;
array2[15574]=30'd231362949;
array2[15575]=30'd231362949;
array2[15576]=30'd231362949;
array2[15577]=30'd231359873;
array2[15578]=30'd231362949;
array2[15579]=30'd231359873;
array2[15580]=30'd234504581;
array2[15581]=30'd231362949;
array2[15582]=30'd231362949;
array2[15583]=30'd230317442;
array2[15584]=30'd229266819;
array2[15585]=30'd231362949;
array2[15586]=30'd231362949;
array2[15587]=30'd231364996;
array2[15588]=30'd231364996;
array2[15589]=30'd231362949;
array2[15590]=30'd229266819;
array2[15591]=30'd231362949;
array2[15592]=30'd231359873;
array2[15593]=30'd231362949;
array2[15594]=30'd231359873;
array2[15595]=30'd231362949;
array2[15596]=30'd229266819;
array2[15597]=30'd231362949;
array2[15598]=30'd229266819;
array2[15599]=30'd231364996;
array2[15600]=30'd231362949;
array2[15601]=30'd231362949;
array2[15602]=30'd229266819;
array2[15603]=30'd231362949;
array2[15604]=30'd234504581;
array2[15605]=30'd231362949;
array2[15606]=30'd227165569;
array2[15607]=30'd231362949;
array2[15608]=30'd231362949;
array2[15609]=30'd231362949;
array2[15610]=30'd231362949;
array2[15611]=30'd229266819;
array2[15612]=30'd231362949;
array2[15613]=30'd230317442;
array2[15614]=30'd230317442;
array2[15615]=30'd231364996;
array2[15616]=30'd231362949;
array2[15617]=30'd231362949;
array2[15618]=30'd231364996;
array2[15619]=30'd228216193;
array2[15620]=30'd231359873;
array2[15621]=30'd231362949;
array2[15622]=30'd230317442;
array2[15623]=30'd231362949;
array2[15624]=30'd230317442;
array2[15625]=30'd230317442;
array2[15626]=30'd231362949;
array2[15627]=30'd230317442;
array2[15628]=30'd231362949;
array2[15629]=30'd228216193;
array2[15630]=30'd231362949;
array2[15631]=30'd231362949;
array2[15632]=30'd231362949;
array2[15633]=30'd230317442;
array2[15634]=30'd230317442;
array2[15635]=30'd231362949;
array2[15636]=30'd231362949;
array2[15637]=30'd229266819;
array2[15638]=30'd234504581;
array2[15639]=30'd228216193;
array2[15640]=30'd231362949;
array2[15641]=30'd231362949;
array2[15642]=30'd231362949;
array2[15643]=30'd231362949;
array2[15644]=30'd231362949;
array2[15645]=30'd234504581;
array2[15646]=30'd231362949;
array2[15647]=30'd231362949;
array2[15648]=30'd212454818;
array2[15649]=30'd231359873;
array2[15650]=30'd227165569;
array2[15651]=30'd231362949;
array2[15652]=30'd234504581;
array2[15653]=30'd228216193;
array2[15654]=30'd231362949;
array2[15655]=30'd229266819;
array2[15656]=30'd231359873;
array2[15657]=30'd231362949;
array2[15658]=30'd231362949;
array2[15659]=30'd231359873;
array2[15660]=30'd231362949;
array2[15661]=30'd231359873;
array2[15662]=30'd231359873;
array2[15663]=30'd231362949;
array2[15664]=30'd229266819;
array2[15665]=30'd230317442;
array2[15666]=30'd225072515;
array2[15667]=30'd228212100;
array2[15668]=30'd229266819;
array2[15669]=30'd231364996;
array2[15670]=30'd229266819;
array2[15671]=30'd231362949;
array2[15672]=30'd229266819;
array2[15673]=30'd231362949;
array2[15674]=30'd234504581;
array2[15675]=30'd231359873;
array2[15676]=30'd227165569;
array2[15677]=30'd231362949;
array2[15678]=30'd231362949;
array2[15679]=30'd228216193;
array2[15680]=30'd231359873;
array2[15681]=30'd231362949;
array2[15682]=30'd231362949;
array2[15683]=30'd231362949;
array2[15684]=30'd229266819;
array2[15685]=30'd231362949;
array2[15686]=30'd231362949;
array2[15687]=30'd229266819;
array2[15688]=30'd231362949;
array2[15689]=30'd231362949;
array2[15690]=30'd229266819;
array2[15691]=30'd229266819;
array2[15692]=30'd229266819;
array2[15693]=30'd231359873;
array2[15694]=30'd231359873;
array2[15695]=30'd231362949;
array2[15696]=30'd229266819;
array2[15697]=30'd231362949;
array2[15698]=30'd228216193;
array2[15699]=30'd228216193;
array2[15700]=30'd231362949;
array2[15701]=30'd231362949;
array2[15702]=30'd231364996;
array2[15703]=30'd230317442;
array2[15704]=30'd231359873;
array2[15705]=30'd231362949;
array2[15706]=30'd231362949;
array2[15707]=30'd234504581;
array2[15708]=30'd231362949;
array2[15709]=30'd230317442;
array2[15710]=30'd231362949;
array2[15711]=30'd229266819;
array2[15712]=30'd231362949;
array2[15713]=30'd231362949;
array2[15714]=30'd231362949;
array2[15715]=30'd231362949;
array2[15716]=30'd229270912;
array2[15717]=30'd229266819;
array2[15718]=30'd230317442;
array2[15719]=30'd231362949;
array2[15720]=30'd231362949;
array2[15721]=30'd231359873;
array2[15722]=30'd231362949;
array2[15723]=30'd231364996;
array2[15724]=30'd231362949;
array2[15725]=30'd231362949;
array2[15726]=30'd231362949;
array2[15727]=30'd231362949;
array2[15728]=30'd231362949;
array2[15729]=30'd231362949;
array2[15730]=30'd231362949;
array2[15731]=30'd231362949;
array2[15732]=30'd231362949;
array2[15733]=30'd231362949;
array2[15734]=30'd234504581;
array2[15735]=30'd229266819;
array2[15736]=30'd231362949;
array2[15737]=30'd229266819;
array2[15738]=30'd231362949;
array2[15739]=30'd234504581;
array2[15740]=30'd234504581;
array2[15741]=30'd229266819;
array2[15742]=30'd231362949;
array2[15743]=30'd228216193;
array2[15744]=30'd212454818;
array2[15745]=30'd234504581;
array2[15746]=30'd227165569;
array2[15747]=30'd231362949;
array2[15748]=30'd231362949;
array2[15749]=30'd229266819;
array2[15750]=30'd229266819;
array2[15751]=30'd231362949;
array2[15752]=30'd229266819;
array2[15753]=30'd231362949;
array2[15754]=30'd231364996;
array2[15755]=30'd231362949;
array2[15756]=30'd231362949;
array2[15757]=30'd229266819;
array2[15758]=30'd231362949;
array2[15759]=30'd228216193;
array2[15760]=30'd229266819;
array2[15761]=30'd231362949;
array2[15762]=30'd195647926;
array2[15763]=30'd319215128;
array2[15764]=30'd260631016;
array2[15765]=30'd212454818;
array2[15766]=30'd186252693;
array2[15767]=30'd228181405;
array2[15768]=30'd231362949;
array2[15769]=30'd228216193;
array2[15770]=30'd229266819;
array2[15771]=30'd231362949;
array2[15772]=30'd231362949;
array2[15773]=30'd231362949;
array2[15774]=30'd231362949;
array2[15775]=30'd227165569;
array2[15776]=30'd231362949;
array2[15777]=30'd231362949;
array2[15778]=30'd231362949;
array2[15779]=30'd230317442;
array2[15780]=30'd231362949;
array2[15781]=30'd229266819;
array2[15782]=30'd231362949;
array2[15783]=30'd231362949;
array2[15784]=30'd231362949;
array2[15785]=30'd230317442;
array2[15786]=30'd229266819;
array2[15787]=30'd228216193;
array2[15788]=30'd231364996;
array2[15789]=30'd231362949;
array2[15790]=30'd231362949;
array2[15791]=30'd231362949;
array2[15792]=30'd231362949;
array2[15793]=30'd231362949;
array2[15794]=30'd229266819;
array2[15795]=30'd229266819;
array2[15796]=30'd234504581;
array2[15797]=30'd231362949;
array2[15798]=30'd230317442;
array2[15799]=30'd231362949;
array2[15800]=30'd231362949;
array2[15801]=30'd228216193;
array2[15802]=30'd231362949;
array2[15803]=30'd230317442;
array2[15804]=30'd230317442;
array2[15805]=30'd229270912;
array2[15806]=30'd229266819;
array2[15807]=30'd231362949;
array2[15808]=30'd229266819;
array2[15809]=30'd231362949;
array2[15810]=30'd234504581;
array2[15811]=30'd231362949;
array2[15812]=30'd231362949;
array2[15813]=30'd231362949;
array2[15814]=30'd229266819;
array2[15815]=30'd230317442;
array2[15816]=30'd231362949;
array2[15817]=30'd231362949;
array2[15818]=30'd229266819;
array2[15819]=30'd231362949;
array2[15820]=30'd231362949;
array2[15821]=30'd231362949;
array2[15822]=30'd231362949;
array2[15823]=30'd229266819;
array2[15824]=30'd231362949;
array2[15825]=30'd231359873;
array2[15826]=30'd227165569;
array2[15827]=30'd231362949;
array2[15828]=30'd231362949;
array2[15829]=30'd230317442;
array2[15830]=30'd229266819;
array2[15831]=30'd229266819;
array2[15832]=30'd229266819;
array2[15833]=30'd234504581;
array2[15834]=30'd231362949;
array2[15835]=30'd229266819;
array2[15836]=30'd231362949;
array2[15837]=30'd234504581;
array2[15838]=30'd238691720;
array2[15839]=30'd234499470;
array2[15840]=30'd212454818;
array2[15841]=30'd234504581;
array2[15842]=30'd227165569;
array2[15843]=30'd231362949;
array2[15844]=30'd231362949;
array2[15845]=30'd231362949;
array2[15846]=30'd231364996;
array2[15847]=30'd231362949;
array2[15848]=30'd231362949;
array2[15849]=30'd231362949;
array2[15850]=30'd234504581;
array2[15851]=30'd229266819;
array2[15852]=30'd231362949;
array2[15853]=30'd229266819;
array2[15854]=30'd231362949;
array2[15855]=30'd231362949;
array2[15856]=30'd231362949;
array2[15857]=30'd229266819;
array2[15858]=30'd195647926;
array2[15859]=30'd645112409;
array2[15860]=30'd566515308;
array2[15861]=30'd538207812;
array2[15862]=30'd538207812;
array2[15863]=30'd383147560;
array2[15864]=30'd207191473;
array2[15865]=30'd193577377;
array2[15866]=30'd207191473;
array2[15867]=30'd234499470;
array2[15868]=30'd231359873;
array2[15869]=30'd231364996;
array2[15870]=30'd229266819;
array2[15871]=30'd231362949;
array2[15872]=30'd231362949;
array2[15873]=30'd231362949;
array2[15874]=30'd231362949;
array2[15875]=30'd231359873;
array2[15876]=30'd227165569;
array2[15877]=30'd231362949;
array2[15878]=30'd234504581;
array2[15879]=30'd231362949;
array2[15880]=30'd231364996;
array2[15881]=30'd229266819;
array2[15882]=30'd229266819;
array2[15883]=30'd229266819;
array2[15884]=30'd231362949;
array2[15885]=30'd231362949;
array2[15886]=30'd228216193;
array2[15887]=30'd231362949;
array2[15888]=30'd231362949;
array2[15889]=30'd229266819;
array2[15890]=30'd230317442;
array2[15891]=30'd231362949;
array2[15892]=30'd229266819;
array2[15893]=30'd230317442;
array2[15894]=30'd231362949;
array2[15895]=30'd231362949;
array2[15896]=30'd231362949;
array2[15897]=30'd231364996;
array2[15898]=30'd231362949;
array2[15899]=30'd229266819;
array2[15900]=30'd230317442;
array2[15901]=30'd231362949;
array2[15902]=30'd231362949;
array2[15903]=30'd231362949;
array2[15904]=30'd229266819;
array2[15905]=30'd231362949;
array2[15906]=30'd231362949;
array2[15907]=30'd229266819;
array2[15908]=30'd229266819;
array2[15909]=30'd231362949;
array2[15910]=30'd230317442;
array2[15911]=30'd231362949;
array2[15912]=30'd229266819;
array2[15913]=30'd231362949;
array2[15914]=30'd229266819;
array2[15915]=30'd230317442;
array2[15916]=30'd231364996;
array2[15917]=30'd234504581;
array2[15918]=30'd231362949;
array2[15919]=30'd231362949;
array2[15920]=30'd231362949;
array2[15921]=30'd228216193;
array2[15922]=30'd230317442;
array2[15923]=30'd231362949;
array2[15924]=30'd231362949;
array2[15925]=30'd229266819;
array2[15926]=30'd231362949;
array2[15927]=30'd231362949;
array2[15928]=30'd231362949;
array2[15929]=30'd231362949;
array2[15930]=30'd229266819;
array2[15931]=30'd231364996;
array2[15932]=30'd228216193;
array2[15933]=30'd616102353;
array2[15934]=30'd777593273;
array2[15935]=30'd281654691;
array2[15936]=30'd212454818;
array2[15937]=30'd234504581;
array2[15938]=30'd228212100;
array2[15939]=30'd234504581;
array2[15940]=30'd234504581;
array2[15941]=30'd231362949;
array2[15942]=30'd231362949;
array2[15943]=30'd231362949;
array2[15944]=30'd231362949;
array2[15945]=30'd231362949;
array2[15946]=30'd234504581;
array2[15947]=30'd231362949;
array2[15948]=30'd231362949;
array2[15949]=30'd229266819;
array2[15950]=30'd231362949;
array2[15951]=30'd229266819;
array2[15952]=30'd229266819;
array2[15953]=30'd231362949;
array2[15954]=30'd207191473;
array2[15955]=30'd645112409;
array2[15956]=30'd858839683;
array2[15957]=30'd865130113;
array2[15958]=30'd858839683;
array2[15959]=30'd727851632;
array2[15960]=30'd565444213;
array2[15961]=30'd645112409;
array2[15962]=30'd506770009;
array2[15963]=30'd195647926;
array2[15964]=30'd195647926;
array2[15965]=30'd212454818;
array2[15966]=30'd228216193;
array2[15967]=30'd230307208;
array2[15968]=30'd228216193;
array2[15969]=30'd229266819;
array2[15970]=30'd229266819;
array2[15971]=30'd231362949;
array2[15972]=30'd231362949;
array2[15973]=30'd234504581;
array2[15974]=30'd234504581;
array2[15975]=30'd227165569;
array2[15976]=30'd231362949;
array2[15977]=30'd231362949;
array2[15978]=30'd231362949;
array2[15979]=30'd230317442;
array2[15980]=30'd231364996;
array2[15981]=30'd231362949;
array2[15982]=30'd231362949;
array2[15983]=30'd231362949;
array2[15984]=30'd231362949;
array2[15985]=30'd228216193;
array2[15986]=30'd229266819;
array2[15987]=30'd234504581;
array2[15988]=30'd231362949;
array2[15989]=30'd229266819;
array2[15990]=30'd231362949;
array2[15991]=30'd229266819;
array2[15992]=30'd231362949;
array2[15993]=30'd231362949;
array2[15994]=30'd228216193;
array2[15995]=30'd229266819;
array2[15996]=30'd231362949;
array2[15997]=30'd230317442;
array2[15998]=30'd231364996;
array2[15999]=30'd230317442;
array2[16000]=30'd228216193;
array2[16001]=30'd231362949;
array2[16002]=30'd231362949;
array2[16003]=30'd231362949;
array2[16004]=30'd228216193;
array2[16005]=30'd231362949;
array2[16006]=30'd231362949;
array2[16007]=30'd234504581;
array2[16008]=30'd229266819;
array2[16009]=30'd231362949;
array2[16010]=30'd231362949;
array2[16011]=30'd231362949;
array2[16012]=30'd231362949;
array2[16013]=30'd231362949;
array2[16014]=30'd231362949;
array2[16015]=30'd234504581;
array2[16016]=30'd231359873;
array2[16017]=30'd231362949;
array2[16018]=30'd231362949;
array2[16019]=30'd229266819;
array2[16020]=30'd229266819;
array2[16021]=30'd231359873;
array2[16022]=30'd231362949;
array2[16023]=30'd231362949;
array2[16024]=30'd231362949;
array2[16025]=30'd229266819;
array2[16026]=30'd231362949;
array2[16027]=30'd231364996;
array2[16028]=30'd221916546;
array2[16029]=30'd719920570;
array2[16030]=30'd970500575;
array2[16031]=30'd281654691;
array2[16032]=30'd212454818;
array2[16033]=30'd234504581;
array2[16034]=30'd227165569;
array2[16035]=30'd231362949;
array2[16036]=30'd234504581;
array2[16037]=30'd231362949;
array2[16038]=30'd231362949;
array2[16039]=30'd231364996;
array2[16040]=30'd231362949;
array2[16041]=30'd231362949;
array2[16042]=30'd228216193;
array2[16043]=30'd228216193;
array2[16044]=30'd230317442;
array2[16045]=30'd230317442;
array2[16046]=30'd229270912;
array2[16047]=30'd229266819;
array2[16048]=30'd231362949;
array2[16049]=30'd230317442;
array2[16050]=30'd221916546;
array2[16051]=30'd319215128;
array2[16052]=30'd805398138;
array2[16053]=30'd858839683;
array2[16054]=30'd865130113;
array2[16055]=30'd865130113;
array2[16056]=30'd865130113;
array2[16057]=30'd865130113;
array2[16058]=30'd828452495;
array2[16059]=30'd727851632;
array2[16060]=30'd727851632;
array2[16061]=30'd483727963;
array2[16062]=30'd190356956;
array2[16063]=30'd190356956;
array2[16064]=30'd213516691;
array2[16065]=30'd225072515;
array2[16066]=30'd227165569;
array2[16067]=30'd228216193;
array2[16068]=30'd231362949;
array2[16069]=30'd231362949;
array2[16070]=30'd229266819;
array2[16071]=30'd230317442;
array2[16072]=30'd231362949;
array2[16073]=30'd228216193;
array2[16074]=30'd231362949;
array2[16075]=30'd230317442;
array2[16076]=30'd231364996;
array2[16077]=30'd231362949;
array2[16078]=30'd231362949;
array2[16079]=30'd231362949;
array2[16080]=30'd231362949;
array2[16081]=30'd231362949;
array2[16082]=30'd231362949;
array2[16083]=30'd230317442;
array2[16084]=30'd234504581;
array2[16085]=30'd229266819;
array2[16086]=30'd229266819;
array2[16087]=30'd231364996;
array2[16088]=30'd234504581;
array2[16089]=30'd231364996;
array2[16090]=30'd231362949;
array2[16091]=30'd230317442;
array2[16092]=30'd231362949;
array2[16093]=30'd228212100;
array2[16094]=30'd231362949;
array2[16095]=30'd231362949;
array2[16096]=30'd234504581;
array2[16097]=30'd229266819;
array2[16098]=30'd231362949;
array2[16099]=30'd228216193;
array2[16100]=30'd230317442;
array2[16101]=30'd229270912;
array2[16102]=30'd229266819;
array2[16103]=30'd231362949;
array2[16104]=30'd229266819;
array2[16105]=30'd231362949;
array2[16106]=30'd231362949;
array2[16107]=30'd231362949;
array2[16108]=30'd231364996;
array2[16109]=30'd231362949;
array2[16110]=30'd229266819;
array2[16111]=30'd230317442;
array2[16112]=30'd231362949;
array2[16113]=30'd234504581;
array2[16114]=30'd229266819;
array2[16115]=30'd231362949;
array2[16116]=30'd231364996;
array2[16117]=30'd228216193;
array2[16118]=30'd225072515;
array2[16119]=30'd231362949;
array2[16120]=30'd231362949;
array2[16121]=30'd234504581;
array2[16122]=30'd231362949;
array2[16123]=30'd231362949;
array2[16124]=30'd227165569;
array2[16125]=30'd464076202;
array2[16126]=30'd616102353;
array2[16127]=30'd262793620;
array2[16128]=30'd212454818;
array2[16129]=30'd234504581;
array2[16130]=30'd227165569;
array2[16131]=30'd231362949;
array2[16132]=30'd234504581;
array2[16133]=30'd231362949;
array2[16134]=30'd231362949;
array2[16135]=30'd230317442;
array2[16136]=30'd231362949;
array2[16137]=30'd231362949;
array2[16138]=30'd228216193;
array2[16139]=30'd229266819;
array2[16140]=30'd231362949;
array2[16141]=30'd230317442;
array2[16142]=30'd230317442;
array2[16143]=30'd231364996;
array2[16144]=30'd228216193;
array2[16145]=30'd231362949;
array2[16146]=30'd231362949;
array2[16147]=30'd195647926;
array2[16148]=30'd764529268;
array2[16149]=30'd865130113;
array2[16150]=30'd865130113;
array2[16151]=30'd858839683;
array2[16152]=30'd865130113;
array2[16153]=30'd858839683;
array2[16154]=30'd858839683;
array2[16155]=30'd858839683;
array2[16156]=30'd858839683;
array2[16157]=30'd805398138;
array2[16158]=30'd764529268;
array2[16159]=30'd677571193;
array2[16160]=30'd347490866;
array2[16161]=30'd190356956;
array2[16162]=30'd260631016;
array2[16163]=30'd221916546;
array2[16164]=30'd225072515;
array2[16165]=30'd231362949;
array2[16166]=30'd231362949;
array2[16167]=30'd231359873;
array2[16168]=30'd231362949;
array2[16169]=30'd231362949;
array2[16170]=30'd231362949;
array2[16171]=30'd231362949;
array2[16172]=30'd228216193;
array2[16173]=30'd228216193;
array2[16174]=30'd231362949;
array2[16175]=30'd231362949;
array2[16176]=30'd229266819;
array2[16177]=30'd231362949;
array2[16178]=30'd230317442;
array2[16179]=30'd229266819;
array2[16180]=30'd234504581;
array2[16181]=30'd228216193;
array2[16182]=30'd231362949;
array2[16183]=30'd231362949;
array2[16184]=30'd231362949;
array2[16185]=30'd231362949;
array2[16186]=30'd231362949;
array2[16187]=30'd231362949;
array2[16188]=30'd230317442;
array2[16189]=30'd230317442;
array2[16190]=30'd231362949;
array2[16191]=30'd231362949;
array2[16192]=30'd231362949;
array2[16193]=30'd229266819;
array2[16194]=30'd231362949;
array2[16195]=30'd230307208;
array2[16196]=30'd231364996;
array2[16197]=30'd231364996;
array2[16198]=30'd231362949;
array2[16199]=30'd230317442;
array2[16200]=30'd229266819;
array2[16201]=30'd231362949;
array2[16202]=30'd231362949;
array2[16203]=30'd231362949;
array2[16204]=30'd231362949;
array2[16205]=30'd231362949;
array2[16206]=30'd227165569;
array2[16207]=30'd231364996;
array2[16208]=30'd229266819;
array2[16209]=30'd229266819;
array2[16210]=30'd229266819;
array2[16211]=30'd228216193;
array2[16212]=30'd231359873;
array2[16213]=30'd231362949;
array2[16214]=30'd229266819;
array2[16215]=30'd231362949;
array2[16216]=30'd231362949;
array2[16217]=30'd603537847;
array2[16218]=30'd777593273;
array2[16219]=30'd719920570;
array2[16220]=30'd304706973;
array2[16221]=30'd532258209;
array2[16222]=30'd719920570;
array2[16223]=30'd262793620;
array2[16224]=30'd212454818;
array2[16225]=30'd234504581;
array2[16226]=30'd227165569;
array2[16227]=30'd231362949;
array2[16228]=30'd234504581;
array2[16229]=30'd231362949;
array2[16230]=30'd231362949;
array2[16231]=30'd229266819;
array2[16232]=30'd231362949;
array2[16233]=30'd228216193;
array2[16234]=30'd231362949;
array2[16235]=30'd234504581;
array2[16236]=30'd231362949;
array2[16237]=30'd231362949;
array2[16238]=30'd231362949;
array2[16239]=30'd231359873;
array2[16240]=30'd228216193;
array2[16241]=30'd231362949;
array2[16242]=30'd231362949;
array2[16243]=30'd195647926;
array2[16244]=30'd764529268;
array2[16245]=30'd865130113;
array2[16246]=30'd865130113;
array2[16247]=30'd865130113;
array2[16248]=30'd858839683;
array2[16249]=30'd858839683;
array2[16250]=30'd858839683;
array2[16251]=30'd858839683;
array2[16252]=30'd858839683;
array2[16253]=30'd858839683;
array2[16254]=30'd865130113;
array2[16255]=30'd851505800;
array2[16256]=30'd805398138;
array2[16257]=30'd790726247;
array2[16258]=30'd631447172;
array2[16259]=30'd319215128;
array2[16260]=30'd212454818;
array2[16261]=30'd234504581;
array2[16262]=30'd234504581;
array2[16263]=30'd229266819;
array2[16264]=30'd231362949;
array2[16265]=30'd231362949;
array2[16266]=30'd231362949;
array2[16267]=30'd231362949;
array2[16268]=30'd234504581;
array2[16269]=30'd231362949;
array2[16270]=30'd231362949;
array2[16271]=30'd231362949;
array2[16272]=30'd229266819;
array2[16273]=30'd231362949;
array2[16274]=30'd229266819;
array2[16275]=30'd231362949;
array2[16276]=30'd234504581;
array2[16277]=30'd231362949;
array2[16278]=30'd229266819;
array2[16279]=30'd231362949;
array2[16280]=30'd231362949;
array2[16281]=30'd231362949;
array2[16282]=30'd231362949;
array2[16283]=30'd234504581;
array2[16284]=30'd231362949;
array2[16285]=30'd231364996;
array2[16286]=30'd229266819;
array2[16287]=30'd231362949;
array2[16288]=30'd231362949;
array2[16289]=30'd234504581;
array2[16290]=30'd231362949;
array2[16291]=30'd227165569;
array2[16292]=30'd231362949;
array2[16293]=30'd231362949;
array2[16294]=30'd231362949;
array2[16295]=30'd229266819;
array2[16296]=30'd231362949;
array2[16297]=30'd228216193;
array2[16298]=30'd231362949;
array2[16299]=30'd231362949;
array2[16300]=30'd231362949;
array2[16301]=30'd231362949;
array2[16302]=30'd231362949;
array2[16303]=30'd234504581;
array2[16304]=30'd231362949;
array2[16305]=30'd231359873;
array2[16306]=30'd231362949;
array2[16307]=30'd231362949;
array2[16308]=30'd231362949;
array2[16309]=30'd229266819;
array2[16310]=30'd231362949;
array2[16311]=30'd234504581;
array2[16312]=30'd234504581;
array2[16313]=30'd532258209;
array2[16314]=30'd670611929;
array2[16315]=30'd670611929;
array2[16316]=30'd304706973;
array2[16317]=30'd464076202;
array2[16318]=30'd670611929;
array2[16319]=30'd262793620;
array2[16320]=30'd212454818;
array2[16321]=30'd234504581;
array2[16322]=30'd234504581;
array2[16323]=30'd230317442;
array2[16324]=30'd229266819;
array2[16325]=30'd229266819;
array2[16326]=30'd231359873;
array2[16327]=30'd231359873;
array2[16328]=30'd227165569;
array2[16329]=30'd234504581;
array2[16330]=30'd234504581;
array2[16331]=30'd228216193;
array2[16332]=30'd231362949;
array2[16333]=30'd231362949;
array2[16334]=30'd229266819;
array2[16335]=30'd231362949;
array2[16336]=30'd230317442;
array2[16337]=30'd231362949;
array2[16338]=30'd231362949;
array2[16339]=30'd195647926;
array2[16340]=30'd764529268;
array2[16341]=30'd851505800;
array2[16342]=30'd865130113;
array2[16343]=30'd865130113;
array2[16344]=30'd858839683;
array2[16345]=30'd858839683;
array2[16346]=30'd858839683;
array2[16347]=30'd858839683;
array2[16348]=30'd858839683;
array2[16349]=30'd858839683;
array2[16350]=30'd858839683;
array2[16351]=30'd858839683;
array2[16352]=30'd858839683;
array2[16353]=30'd858839683;
array2[16354]=30'd828452495;
array2[16355]=30'd566515308;
array2[16356]=30'd186252693;
array2[16357]=30'd230317442;
array2[16358]=30'd231364996;
array2[16359]=30'd229266819;
array2[16360]=30'd230317442;
array2[16361]=30'd231362949;
array2[16362]=30'd231364996;
array2[16363]=30'd228216193;
array2[16364]=30'd228216193;
array2[16365]=30'd231362949;
array2[16366]=30'd231362949;
array2[16367]=30'd230317442;
array2[16368]=30'd230317442;
array2[16369]=30'd229266819;
array2[16370]=30'd231362949;
array2[16371]=30'd229266819;
array2[16372]=30'd231362949;
array2[16373]=30'd228216193;
array2[16374]=30'd229266819;
array2[16375]=30'd231362949;
array2[16376]=30'd230317442;
array2[16377]=30'd230317442;
array2[16378]=30'd231364996;
array2[16379]=30'd231362949;
array2[16380]=30'd231362949;
array2[16381]=30'd231362949;
array2[16382]=30'd231362949;
array2[16383]=30'd231362949;
array2[16384]=30'd227165569;
array2[16385]=30'd231362949;
array2[16386]=30'd231362949;
array2[16387]=30'd231364996;
array2[16388]=30'd230317442;
array2[16389]=30'd230317442;
array2[16390]=30'd228216193;
array2[16391]=30'd231359873;
array2[16392]=30'd231362949;
array2[16393]=30'd230317442;
array2[16394]=30'd231362949;
array2[16395]=30'd231362949;
array2[16396]=30'd231362949;
array2[16397]=30'd230317442;
array2[16398]=30'd229266819;
array2[16399]=30'd234504581;
array2[16400]=30'd228216193;
array2[16401]=30'd231362949;
array2[16402]=30'd231362949;
array2[16403]=30'd229266819;
array2[16404]=30'd231362949;
array2[16405]=30'd231362949;
array2[16406]=30'd234504581;
array2[16407]=30'd231362949;
array2[16408]=30'd231362949;
array2[16409]=30'd229266819;
array2[16410]=30'd228212100;
array2[16411]=30'd221916546;
array2[16412]=30'd231362949;
array2[16413]=30'd425297329;
array2[16414]=30'd616102353;
array2[16415]=30'd262793620;
array2[16416]=30'd228181405;
array2[16417]=30'd234504581;
array2[16418]=30'd227159434;
array2[16419]=30'd228216193;
array2[16420]=30'd231364996;
array2[16421]=30'd229266819;
array2[16422]=30'd229266819;
array2[16423]=30'd231362949;
array2[16424]=30'd231364996;
array2[16425]=30'd231362949;
array2[16426]=30'd227165569;
array2[16427]=30'd231362949;
array2[16428]=30'd231362949;
array2[16429]=30'd230317442;
array2[16430]=30'd231362949;
array2[16431]=30'd231364996;
array2[16432]=30'd230317442;
array2[16433]=30'd231364996;
array2[16434]=30'd231364996;
array2[16435]=30'd207191473;
array2[16436]=30'd565444213;
array2[16437]=30'd819020415;
array2[16438]=30'd858839683;
array2[16439]=30'd858839683;
array2[16440]=30'd858839683;
array2[16441]=30'd858839683;
array2[16442]=30'd858839683;
array2[16443]=30'd858839683;
array2[16444]=30'd858839683;
array2[16445]=30'd858839683;
array2[16446]=30'd858839683;
array2[16447]=30'd858839683;
array2[16448]=30'd858839683;
array2[16449]=30'd858839683;
array2[16450]=30'd805398138;
array2[16451]=30'd450208341;
array2[16452]=30'd212454818;
array2[16453]=30'd231362949;
array2[16454]=30'd231362949;
array2[16455]=30'd231362949;
array2[16456]=30'd231362949;
array2[16457]=30'd229266819;
array2[16458]=30'd231364996;
array2[16459]=30'd231362949;
array2[16460]=30'd228216193;
array2[16461]=30'd228216193;
array2[16462]=30'd231362949;
array2[16463]=30'd230317442;
array2[16464]=30'd230317442;
array2[16465]=30'd230317442;
array2[16466]=30'd231362949;
array2[16467]=30'd231362949;
array2[16468]=30'd231362949;
array2[16469]=30'd231362949;
array2[16470]=30'd228216193;
array2[16471]=30'd231362949;
array2[16472]=30'd231362949;
array2[16473]=30'd231364996;
array2[16474]=30'd231362949;
array2[16475]=30'd229266819;
array2[16476]=30'd231362949;
array2[16477]=30'd231362949;
array2[16478]=30'd231362949;
array2[16479]=30'd231362949;
array2[16480]=30'd231364996;
array2[16481]=30'd227165569;
array2[16482]=30'd231364996;
array2[16483]=30'd230317442;
array2[16484]=30'd230317442;
array2[16485]=30'd231362949;
array2[16486]=30'd231362949;
array2[16487]=30'd229266819;
array2[16488]=30'd228216193;
array2[16489]=30'd231362949;
array2[16490]=30'd231362949;
array2[16491]=30'd231362949;
array2[16492]=30'd230317442;
array2[16493]=30'd230317442;
array2[16494]=30'd231362949;
array2[16495]=30'd231362949;
array2[16496]=30'd229266819;
array2[16497]=30'd234504581;
array2[16498]=30'd231362949;
array2[16499]=30'd231362949;
array2[16500]=30'd227165569;
array2[16501]=30'd229266819;
array2[16502]=30'd231362949;
array2[16503]=30'd231362949;
array2[16504]=30'd231362949;
array2[16505]=30'd229266819;
array2[16506]=30'd231362949;
array2[16507]=30'd231364996;
array2[16508]=30'd231362949;
array2[16509]=30'd664345022;
array2[16510]=30'd970500575;
array2[16511]=30'd281654691;
array2[16512]=30'd228181405;
array2[16513]=30'd234504581;
array2[16514]=30'd234504581;
array2[16515]=30'd231362949;
array2[16516]=30'd231362949;
array2[16517]=30'd229266819;
array2[16518]=30'd231362949;
array2[16519]=30'd231362949;
array2[16520]=30'd231359873;
array2[16521]=30'd234504581;
array2[16522]=30'd234504581;
array2[16523]=30'd234504581;
array2[16524]=30'd231362949;
array2[16525]=30'd231362949;
array2[16526]=30'd229266819;
array2[16527]=30'd229266819;
array2[16528]=30'd229266819;
array2[16529]=30'd230317442;
array2[16530]=30'd231364996;
array2[16531]=30'd227159434;
array2[16532]=30'd281508345;
array2[16533]=30'd805398138;
array2[16534]=30'd858839683;
array2[16535]=30'd858839683;
array2[16536]=30'd858839683;
array2[16537]=30'd858839683;
array2[16538]=30'd858839683;
array2[16539]=30'd858839683;
array2[16540]=30'd858839683;
array2[16541]=30'd858839683;
array2[16542]=30'd858839683;
array2[16543]=30'd865130113;
array2[16544]=30'd865130113;
array2[16545]=30'd858839683;
array2[16546]=30'd708987491;
array2[16547]=30'd195647926;
array2[16548]=30'd229270912;
array2[16549]=30'd231362949;
array2[16550]=30'd231362949;
array2[16551]=30'd229266819;
array2[16552]=30'd231362949;
array2[16553]=30'd231362949;
array2[16554]=30'd231362949;
array2[16555]=30'd231359873;
array2[16556]=30'd238691720;
array2[16557]=30'd231362949;
array2[16558]=30'd231362949;
array2[16559]=30'd229266819;
array2[16560]=30'd229266819;
array2[16561]=30'd231362949;
array2[16562]=30'd230317442;
array2[16563]=30'd231362949;
array2[16564]=30'd231364996;
array2[16565]=30'd229266819;
array2[16566]=30'd229266819;
array2[16567]=30'd228216193;
array2[16568]=30'd231362949;
array2[16569]=30'd234504581;
array2[16570]=30'd234504581;
array2[16571]=30'd234504581;
array2[16572]=30'd231362949;
array2[16573]=30'd231362949;
array2[16574]=30'd228216193;
array2[16575]=30'd231362949;
array2[16576]=30'd231362949;
array2[16577]=30'd229266819;
array2[16578]=30'd231362949;
array2[16579]=30'd231362949;
array2[16580]=30'd231359873;
array2[16581]=30'd231362949;
array2[16582]=30'd231359873;
array2[16583]=30'd231362949;
array2[16584]=30'd231362949;
array2[16585]=30'd231362949;
array2[16586]=30'd231362949;
array2[16587]=30'd231359873;
array2[16588]=30'd231362949;
array2[16589]=30'd229266819;
array2[16590]=30'd229266819;
array2[16591]=30'd231362949;
array2[16592]=30'd231362949;
array2[16593]=30'd234504581;
array2[16594]=30'd231364996;
array2[16595]=30'd231362949;
array2[16596]=30'd228216193;
array2[16597]=30'd231362949;
array2[16598]=30'd234504581;
array2[16599]=30'd231362949;
array2[16600]=30'd231362949;
array2[16601]=30'd231362949;
array2[16602]=30'd229266819;
array2[16603]=30'd231362949;
array2[16604]=30'd231359873;
array2[16605]=30'd472496545;
array2[16606]=30'd664345022;
array2[16607]=30'd256519562;
array2[16608]=30'd212454818;
array2[16609]=30'd234504581;
array2[16610]=30'd228212100;
array2[16611]=30'd229266819;
array2[16612]=30'd231364996;
array2[16613]=30'd230317442;
array2[16614]=30'd229266819;
array2[16615]=30'd229266819;
array2[16616]=30'd231362949;
array2[16617]=30'd234504581;
array2[16618]=30'd234504581;
array2[16619]=30'd227165569;
array2[16620]=30'd231362949;
array2[16621]=30'd231362949;
array2[16622]=30'd231362949;
array2[16623]=30'd231362949;
array2[16624]=30'd231359873;
array2[16625]=30'd231362949;
array2[16626]=30'd231359873;
array2[16627]=30'd227159434;
array2[16628]=30'd249001484;
array2[16629]=30'd764529268;
array2[16630]=30'd851505800;
array2[16631]=30'd858839683;
array2[16632]=30'd851505800;
array2[16633]=30'd851505800;
array2[16634]=30'd851505800;
array2[16635]=30'd858839683;
array2[16636]=30'd851505800;
array2[16637]=30'd851505800;
array2[16638]=30'd851505800;
array2[16639]=30'd858839683;
array2[16640]=30'd865130113;
array2[16641]=30'd851505800;
array2[16642]=30'd646130287;
array2[16643]=30'd179916222;
array2[16644]=30'd228216193;
array2[16645]=30'd231359873;
array2[16646]=30'd229266819;
array2[16647]=30'd229266819;
array2[16648]=30'd231359873;
array2[16649]=30'd231359873;
array2[16650]=30'd231362949;
array2[16651]=30'd231362949;
array2[16652]=30'd234504581;
array2[16653]=30'd227165569;
array2[16654]=30'd228216193;
array2[16655]=30'd231362949;
array2[16656]=30'd231362949;
array2[16657]=30'd234504581;
array2[16658]=30'd231359873;
array2[16659]=30'd231362949;
array2[16660]=30'd231362949;
array2[16661]=30'd231362949;
array2[16662]=30'd231362949;
array2[16663]=30'd234504581;
array2[16664]=30'd231362949;
array2[16665]=30'd234504581;
array2[16666]=30'd231362949;
array2[16667]=30'd229266819;
array2[16668]=30'd229266819;
array2[16669]=30'd230317442;
array2[16670]=30'd229266819;
array2[16671]=30'd234504581;
array2[16672]=30'd231362949;
array2[16673]=30'd229266819;
array2[16674]=30'd231362949;
array2[16675]=30'd231362949;
array2[16676]=30'd231362949;
array2[16677]=30'd231362949;
array2[16678]=30'd231362949;
array2[16679]=30'd229266819;
array2[16680]=30'd231362949;
array2[16681]=30'd231362949;
array2[16682]=30'd231364996;
array2[16683]=30'd230317442;
array2[16684]=30'd230317442;
array2[16685]=30'd231362949;
array2[16686]=30'd229266819;
array2[16687]=30'd231362949;
array2[16688]=30'd229266819;
array2[16689]=30'd231362949;
array2[16690]=30'd231362949;
array2[16691]=30'd230317442;
array2[16692]=30'd231362949;
array2[16693]=30'd229266819;
array2[16694]=30'd231362949;
array2[16695]=30'd231362949;
array2[16696]=30'd231362949;
array2[16697]=30'd229266819;
array2[16698]=30'd231362949;
array2[16699]=30'd231362949;
array2[16700]=30'd229270912;
array2[16701]=30'd231362949;
array2[16702]=30'd234504581;
array2[16703]=30'd228216193;
array2[16704]=30'd212454818;
array2[16705]=30'd234504581;
array2[16706]=30'd227165569;
array2[16707]=30'd231362949;
array2[16708]=30'd234504581;
array2[16709]=30'd231362949;
array2[16710]=30'd231362949;
array2[16711]=30'd230317442;
array2[16712]=30'd231362949;
array2[16713]=30'd234504581;
array2[16714]=30'd228216193;
array2[16715]=30'd231362949;
array2[16716]=30'd231362949;
array2[16717]=30'd228216193;
array2[16718]=30'd228216193;
array2[16719]=30'd231364996;
array2[16720]=30'd231362949;
array2[16721]=30'd231364996;
array2[16722]=30'd231362949;
array2[16723]=30'd234504581;
array2[16724]=30'd213516691;
array2[16725]=30'd281508345;
array2[16726]=30'd281508345;
array2[16727]=30'd281508345;
array2[16728]=30'd281508345;
array2[16729]=30'd281508345;
array2[16730]=30'd265736724;
array2[16731]=30'd281508345;
array2[16732]=30'd281508345;
array2[16733]=30'd265736724;
array2[16734]=30'd265736724;
array2[16735]=30'd319215128;
array2[16736]=30'd764529268;
array2[16737]=30'd764529268;
array2[16738]=30'd281508345;
array2[16739]=30'd228181405;
array2[16740]=30'd225072515;
array2[16741]=30'd236604812;
array2[16742]=30'd234504581;
array2[16743]=30'd225072515;
array2[16744]=30'd228216193;
array2[16745]=30'd231359873;
array2[16746]=30'd229266819;
array2[16747]=30'd229266819;
array2[16748]=30'd231362949;
array2[16749]=30'd229266819;
array2[16750]=30'd231362949;
array2[16751]=30'd231362949;
array2[16752]=30'd228216193;
array2[16753]=30'd234504581;
array2[16754]=30'd228216193;
array2[16755]=30'd231364996;
array2[16756]=30'd231362949;
array2[16757]=30'd229266819;
array2[16758]=30'd230317442;
array2[16759]=30'd231362949;
array2[16760]=30'd231359873;
array2[16761]=30'd231362949;
array2[16762]=30'd231362949;
array2[16763]=30'd230317442;
array2[16764]=30'd231364996;
array2[16765]=30'd228212100;
array2[16766]=30'd231364996;
array2[16767]=30'd230317442;
array2[16768]=30'd231362949;
array2[16769]=30'd228216193;
array2[16770]=30'd231364996;
array2[16771]=30'd231362949;
array2[16772]=30'd231362949;
array2[16773]=30'd229266819;
array2[16774]=30'd231364996;
array2[16775]=30'd231362949;
array2[16776]=30'd230317442;
array2[16777]=30'd230317442;
array2[16778]=30'd231362949;
array2[16779]=30'd231364996;
array2[16780]=30'd227165569;
array2[16781]=30'd228216193;
array2[16782]=30'd231362949;
array2[16783]=30'd231364996;
array2[16784]=30'd231362949;
array2[16785]=30'd231362949;
array2[16786]=30'd230317442;
array2[16787]=30'd230317442;
array2[16788]=30'd231362949;
array2[16789]=30'd228216193;
array2[16790]=30'd231359873;
array2[16791]=30'd231364996;
array2[16792]=30'd231364996;
array2[16793]=30'd228216193;
array2[16794]=30'd229266819;
array2[16795]=30'd231362949;
array2[16796]=30'd230317442;
array2[16797]=30'd229266819;
array2[16798]=30'd231359873;
array2[16799]=30'd228216193;
array2[16800]=30'd212454818;
array2[16801]=30'd234504581;
array2[16802]=30'd227165569;
array2[16803]=30'd231362949;
array2[16804]=30'd234504581;
array2[16805]=30'd231362949;
array2[16806]=30'd231362949;
array2[16807]=30'd230317442;
array2[16808]=30'd231362949;
array2[16809]=30'd234504581;
array2[16810]=30'd230317442;
array2[16811]=30'd230317442;
array2[16812]=30'd231364996;
array2[16813]=30'd229266819;
array2[16814]=30'd228216193;
array2[16815]=30'd231362949;
array2[16816]=30'd231362949;
array2[16817]=30'd231362949;
array2[16818]=30'd231362949;
array2[16819]=30'd234504581;
array2[16820]=30'd231362949;
array2[16821]=30'd229266819;
array2[16822]=30'd228216193;
array2[16823]=30'd227165569;
array2[16824]=30'd229266819;
array2[16825]=30'd228216193;
array2[16826]=30'd230307208;
array2[16827]=30'd230307208;
array2[16828]=30'd227165569;
array2[16829]=30'd230307208;
array2[16830]=30'd227159434;
array2[16831]=30'd190356956;
array2[16832]=30'd790726247;
array2[16833]=30'd764529268;
array2[16834]=30'd249001484;
array2[16835]=30'd249001484;
array2[16836]=30'd249001484;
array2[16837]=30'd249001484;
array2[16838]=30'd249001484;
array2[16839]=30'd179916222;
array2[16840]=30'd231362949;
array2[16841]=30'd231362949;
array2[16842]=30'd231362949;
array2[16843]=30'd231359873;
array2[16844]=30'd231362949;
array2[16845]=30'd231362949;
array2[16846]=30'd230317442;
array2[16847]=30'd231364996;
array2[16848]=30'd231362949;
array2[16849]=30'd231362949;
array2[16850]=30'd231362949;
array2[16851]=30'd229266819;
array2[16852]=30'd231362949;
array2[16853]=30'd231362949;
array2[16854]=30'd230317442;
array2[16855]=30'd234504581;
array2[16856]=30'd231362949;
array2[16857]=30'd230317442;
array2[16858]=30'd230317442;
array2[16859]=30'd228216193;
array2[16860]=30'd229266819;
array2[16861]=30'd231362949;
array2[16862]=30'd231364996;
array2[16863]=30'd231362949;
array2[16864]=30'd228212100;
array2[16865]=30'd231362949;
array2[16866]=30'd230317442;
array2[16867]=30'd231362949;
array2[16868]=30'd231362949;
array2[16869]=30'd231359873;
array2[16870]=30'd231364996;
array2[16871]=30'd231362949;
array2[16872]=30'd231362949;
array2[16873]=30'd228216193;
array2[16874]=30'd234504581;
array2[16875]=30'd231362949;
array2[16876]=30'd231362949;
array2[16877]=30'd230317442;
array2[16878]=30'd229266819;
array2[16879]=30'd231362949;
array2[16880]=30'd230317442;
array2[16881]=30'd231362949;
array2[16882]=30'd234504581;
array2[16883]=30'd231362949;
array2[16884]=30'd231364996;
array2[16885]=30'd234504581;
array2[16886]=30'd229266819;
array2[16887]=30'd231362949;
array2[16888]=30'd231362949;
array2[16889]=30'd231359873;
array2[16890]=30'd229266819;
array2[16891]=30'd234504581;
array2[16892]=30'd230317442;
array2[16893]=30'd234504581;
array2[16894]=30'd230307208;
array2[16895]=30'd230317442;
array2[16896]=30'd212454818;
array2[16897]=30'd234504581;
array2[16898]=30'd227165569;
array2[16899]=30'd231364996;
array2[16900]=30'd231362949;
array2[16901]=30'd229266819;
array2[16902]=30'd231362949;
array2[16903]=30'd230317442;
array2[16904]=30'd234504581;
array2[16905]=30'd234504581;
array2[16906]=30'd234504581;
array2[16907]=30'd231362949;
array2[16908]=30'd231362949;
array2[16909]=30'd231362949;
array2[16910]=30'd229266819;
array2[16911]=30'd231362949;
array2[16912]=30'd229266819;
array2[16913]=30'd231359873;
array2[16914]=30'd231362949;
array2[16915]=30'd228216193;
array2[16916]=30'd228216193;
array2[16917]=30'd231364996;
array2[16918]=30'd231364996;
array2[16919]=30'd231362949;
array2[16920]=30'd228216193;
array2[16921]=30'd231362949;
array2[16922]=30'd231359873;
array2[16923]=30'd228216193;
array2[16924]=30'd231362949;
array2[16925]=30'd231362949;
array2[16926]=30'd213516691;
array2[16927]=30'd383147560;
array2[16928]=30'd790726247;
array2[16929]=30'd865130113;
array2[16930]=30'd858839683;
array2[16931]=30'd851505800;
array2[16932]=30'd858839683;
array2[16933]=30'd819020415;
array2[16934]=30'd645112409;
array2[16935]=30'd260631016;
array2[16936]=30'd234504581;
array2[16937]=30'd228212100;
array2[16938]=30'd229266819;
array2[16939]=30'd231364996;
array2[16940]=30'd231362949;
array2[16941]=30'd231362949;
array2[16942]=30'd231362949;
array2[16943]=30'd231359873;
array2[16944]=30'd231362949;
array2[16945]=30'd229266819;
array2[16946]=30'd231364996;
array2[16947]=30'd230317442;
array2[16948]=30'd231362949;
array2[16949]=30'd230317442;
array2[16950]=30'd229266819;
array2[16951]=30'd234504581;
array2[16952]=30'd231362949;
array2[16953]=30'd229266819;
array2[16954]=30'd231362949;
array2[16955]=30'd229266819;
array2[16956]=30'd231362949;
array2[16957]=30'd231364996;
array2[16958]=30'd234504581;
array2[16959]=30'd229266819;
array2[16960]=30'd231362949;
array2[16961]=30'd231362949;
array2[16962]=30'd231362949;
array2[16963]=30'd230307208;
array2[16964]=30'd230317442;
array2[16965]=30'd229266819;
array2[16966]=30'd230317442;
array2[16967]=30'd231362949;
array2[16968]=30'd230317442;
array2[16969]=30'd231364996;
array2[16970]=30'd231362949;
array2[16971]=30'd228216193;
array2[16972]=30'd231359873;
array2[16973]=30'd231364996;
array2[16974]=30'd229266819;
array2[16975]=30'd229266819;
array2[16976]=30'd231362949;
array2[16977]=30'd227165569;
array2[16978]=30'd231362949;
array2[16979]=30'd234504581;
array2[16980]=30'd234504581;
array2[16981]=30'd231362949;
array2[16982]=30'd234504581;
array2[16983]=30'd228216193;
array2[16984]=30'd231362949;
array2[16985]=30'd231362949;
array2[16986]=30'd231362949;
array2[16987]=30'd231362949;
array2[16988]=30'd231364996;
array2[16989]=30'd234504581;
array2[16990]=30'd228216193;
array2[16991]=30'd231359873;
array2[16992]=30'd212454818;
array2[16993]=30'd231359873;
array2[16994]=30'd229266819;
array2[16995]=30'd229266819;
array2[16996]=30'd231362949;
array2[16997]=30'd231362949;
array2[16998]=30'd231362949;
array2[16999]=30'd231362949;
array2[17000]=30'd231359873;
array2[17001]=30'd227165569;
array2[17002]=30'd231362949;
array2[17003]=30'd231362949;
array2[17004]=30'd231362949;
array2[17005]=30'd231364996;
array2[17006]=30'd231362949;
array2[17007]=30'd229266819;
array2[17008]=30'd231359873;
array2[17009]=30'd231362949;
array2[17010]=30'd231362949;
array2[17011]=30'd229266819;
array2[17012]=30'd231362949;
array2[17013]=30'd231362949;
array2[17014]=30'd231362949;
array2[17015]=30'd229266819;
array2[17016]=30'd229266819;
array2[17017]=30'd231362949;
array2[17018]=30'd231364996;
array2[17019]=30'd231362949;
array2[17020]=30'd231362949;
array2[17021]=30'd231362949;
array2[17022]=30'd207191473;
array2[17023]=30'd631447172;
array2[17024]=30'd828452495;
array2[17025]=30'd805398138;
array2[17026]=30'd645112409;
array2[17027]=30'd645112409;
array2[17028]=30'd764529268;
array2[17029]=30'd823228019;
array2[17030]=30'd319215128;
array2[17031]=30'd225072515;
array2[17032]=30'd231364996;
array2[17033]=30'd231364996;
array2[17034]=30'd230317442;
array2[17035]=30'd229266819;
array2[17036]=30'd231362949;
array2[17037]=30'd231359873;
array2[17038]=30'd231362949;
array2[17039]=30'd229266819;
array2[17040]=30'd231362949;
array2[17041]=30'd230317442;
array2[17042]=30'd231362949;
array2[17043]=30'd230317442;
array2[17044]=30'd231362949;
array2[17045]=30'd231362949;
array2[17046]=30'd231362949;
array2[17047]=30'd231364996;
array2[17048]=30'd231362949;
array2[17049]=30'd229266819;
array2[17050]=30'd229266819;
array2[17051]=30'd231362949;
array2[17052]=30'd231362949;
array2[17053]=30'd230317442;
array2[17054]=30'd231364996;
array2[17055]=30'd230317442;
array2[17056]=30'd231362949;
array2[17057]=30'd227165569;
array2[17058]=30'd230317442;
array2[17059]=30'd231362949;
array2[17060]=30'd231362949;
array2[17061]=30'd231364996;
array2[17062]=30'd228216193;
array2[17063]=30'd229266819;
array2[17064]=30'd230317442;
array2[17065]=30'd231364996;
array2[17066]=30'd231362949;
array2[17067]=30'd229266819;
array2[17068]=30'd231362949;
array2[17069]=30'd230317442;
array2[17070]=30'd231362949;
array2[17071]=30'd228212100;
array2[17072]=30'd231362949;
array2[17073]=30'd231362949;
array2[17074]=30'd230317442;
array2[17075]=30'd230317442;
array2[17076]=30'd228216193;
array2[17077]=30'd231362949;
array2[17078]=30'd231362949;
array2[17079]=30'd231364996;
array2[17080]=30'd229266819;
array2[17081]=30'd230317442;
array2[17082]=30'd231362949;
array2[17083]=30'd231362949;
array2[17084]=30'd231364996;
array2[17085]=30'd231362949;
array2[17086]=30'd231362949;
array2[17087]=30'd227165569;
array2[17088]=30'd212454818;
array2[17089]=30'd234504581;
array2[17090]=30'd227165569;
array2[17091]=30'd231362949;
array2[17092]=30'd231362949;
array2[17093]=30'd229266819;
array2[17094]=30'd231362949;
array2[17095]=30'd231362949;
array2[17096]=30'd231362949;
array2[17097]=30'd234504581;
array2[17098]=30'd229266819;
array2[17099]=30'd231359873;
array2[17100]=30'd231362949;
array2[17101]=30'd228216193;
array2[17102]=30'd229266819;
array2[17103]=30'd231362949;
array2[17104]=30'd231362949;
array2[17105]=30'd231362949;
array2[17106]=30'd231362949;
array2[17107]=30'd231362949;
array2[17108]=30'd231362949;
array2[17109]=30'd231362949;
array2[17110]=30'd231362949;
array2[17111]=30'd231362949;
array2[17112]=30'd229266819;
array2[17113]=30'd231362949;
array2[17114]=30'd229266819;
array2[17115]=30'd234504581;
array2[17116]=30'd231362949;
array2[17117]=30'd229266819;
array2[17118]=30'd207191473;
array2[17119]=30'd450208341;
array2[17120]=30'd566515308;
array2[17121]=30'd483727963;
array2[17122]=30'd207191473;
array2[17123]=30'd179916222;
array2[17124]=30'd506770009;
array2[17125]=30'd645112409;
array2[17126]=30'd249001484;
array2[17127]=30'd221916546;
array2[17128]=30'd225072515;
array2[17129]=30'd225072515;
array2[17130]=30'd228216193;
array2[17131]=30'd231362949;
array2[17132]=30'd231362949;
array2[17133]=30'd234504581;
array2[17134]=30'd234504581;
array2[17135]=30'd227165569;
array2[17136]=30'd231362949;
array2[17137]=30'd231362949;
array2[17138]=30'd229266819;
array2[17139]=30'd230317442;
array2[17140]=30'd231362949;
array2[17141]=30'd231362949;
array2[17142]=30'd231362949;
array2[17143]=30'd230317442;
array2[17144]=30'd228216193;
array2[17145]=30'd225072515;
array2[17146]=30'd225072515;
array2[17147]=30'd227165569;
array2[17148]=30'd234504581;
array2[17149]=30'd231362949;
array2[17150]=30'd229266819;
array2[17151]=30'd231362949;
array2[17152]=30'd228216193;
array2[17153]=30'd234504581;
array2[17154]=30'd230317442;
array2[17155]=30'd231362949;
array2[17156]=30'd229266819;
array2[17157]=30'd231362949;
array2[17158]=30'd231362949;
array2[17159]=30'd231362949;
array2[17160]=30'd231362949;
array2[17161]=30'd229266819;
array2[17162]=30'd231364996;
array2[17163]=30'd229266819;
array2[17164]=30'd229266819;
array2[17165]=30'd231362949;
array2[17166]=30'd231362949;
array2[17167]=30'd231359873;
array2[17168]=30'd231362949;
array2[17169]=30'd227165569;
array2[17170]=30'd231362949;
array2[17171]=30'd231362949;
array2[17172]=30'd231362949;
array2[17173]=30'd231362949;
array2[17174]=30'd229266819;
array2[17175]=30'd231362949;
array2[17176]=30'd231362949;
array2[17177]=30'd231362949;
array2[17178]=30'd231362949;
array2[17179]=30'd228216193;
array2[17180]=30'd229266819;
array2[17181]=30'd231362949;
array2[17182]=30'd231362949;
array2[17183]=30'd229266819;
array2[17184]=30'd212454818;
array2[17185]=30'd377085336;
array2[17186]=30'd425297329;
array2[17187]=30'd227159434;
array2[17188]=30'd227165569;
array2[17189]=30'd229266819;
array2[17190]=30'd229266819;
array2[17191]=30'd231359873;
array2[17192]=30'd231359873;
array2[17193]=30'd231362949;
array2[17194]=30'd231362949;
array2[17195]=30'd231362949;
array2[17196]=30'd227165569;
array2[17197]=30'd231362949;
array2[17198]=30'd231362949;
array2[17199]=30'd231362949;
array2[17200]=30'd231362949;
array2[17201]=30'd228216193;
array2[17202]=30'd231362949;
array2[17203]=30'd231362949;
array2[17204]=30'd229266819;
array2[17205]=30'd228216193;
array2[17206]=30'd231362949;
array2[17207]=30'd231362949;
array2[17208]=30'd338288022;
array2[17209]=30'd464076202;
array2[17210]=30'd238691720;
array2[17211]=30'd227165569;
array2[17212]=30'd234504581;
array2[17213]=30'd231362949;
array2[17214]=30'd220861839;
array2[17215]=30'd213516691;
array2[17216]=30'd213516691;
array2[17217]=30'd213516691;
array2[17218]=30'd234504581;
array2[17219]=30'd212454818;
array2[17220]=30'd295074390;
array2[17221]=30'd357913199;
array2[17222]=30'd178773498;
array2[17223]=30'd150539724;
array2[17224]=30'd150539724;
array2[17225]=30'd150539724;
array2[17226]=30'd193577377;
array2[17227]=30'd231362949;
array2[17228]=30'd231362949;
array2[17229]=30'd234504581;
array2[17230]=30'd231362949;
array2[17231]=30'd231362949;
array2[17232]=30'd231362949;
array2[17233]=30'd231362949;
array2[17234]=30'd231362949;
array2[17235]=30'd234504581;
array2[17236]=30'd234504581;
array2[17237]=30'd231362949;
array2[17238]=30'd231362949;
array2[17239]=30'd229266819;
array2[17240]=30'd195647926;
array2[17241]=30'd179916222;
array2[17242]=30'd179916222;
array2[17243]=30'd207191473;
array2[17244]=30'd221916546;
array2[17245]=30'd221916546;
array2[17246]=30'd227165569;
array2[17247]=30'd231362949;
array2[17248]=30'd234504581;
array2[17249]=30'd231362949;
array2[17250]=30'd231362949;
array2[17251]=30'd231362949;
array2[17252]=30'd231362949;
array2[17253]=30'd231362949;
array2[17254]=30'd231359873;
array2[17255]=30'd231362949;
array2[17256]=30'd231362949;
array2[17257]=30'd231362949;
array2[17258]=30'd230317442;
array2[17259]=30'd229266819;
array2[17260]=30'd231362949;
array2[17261]=30'd230317442;
array2[17262]=30'd231362949;
array2[17263]=30'd228216193;
array2[17264]=30'd229266819;
array2[17265]=30'd231362949;
array2[17266]=30'd231362949;
array2[17267]=30'd231362949;
array2[17268]=30'd231364996;
array2[17269]=30'd234504581;
array2[17270]=30'd229266819;
array2[17271]=30'd231362949;
array2[17272]=30'd231362949;
array2[17273]=30'd231362949;
array2[17274]=30'd231362949;
array2[17275]=30'd231362949;
array2[17276]=30'd231362949;
array2[17277]=30'd231362949;
array2[17278]=30'd229266819;
array2[17279]=30'd231362949;
array2[17280]=30'd338288022;
array2[17281]=30'd664345022;
array2[17282]=30'd777593273;
array2[17283]=30'd377085336;
array2[17284]=30'd256519562;
array2[17285]=30'd229270912;
array2[17286]=30'd229270912;
array2[17287]=30'd231362949;
array2[17288]=30'd229266819;
array2[17289]=30'd231362949;
array2[17290]=30'd229266819;
array2[17291]=30'd229266819;
array2[17292]=30'd231362949;
array2[17293]=30'd231362949;
array2[17294]=30'd230317442;
array2[17295]=30'd230317442;
array2[17296]=30'd231362949;
array2[17297]=30'd228216193;
array2[17298]=30'd230317442;
array2[17299]=30'd231362949;
array2[17300]=30'd234504581;
array2[17301]=30'd229266819;
array2[17302]=30'd231362949;
array2[17303]=30'd227165569;
array2[17304]=30'd532258209;
array2[17305]=30'd822672828;
array2[17306]=30'd425297329;
array2[17307]=30'd256519562;
array2[17308]=30'd229270912;
array2[17309]=30'd230317442;
array2[17310]=30'd231362949;
array2[17311]=30'd231362949;
array2[17312]=30'd231362949;
array2[17313]=30'd231362949;
array2[17314]=30'd231362949;
array2[17315]=30'd186252693;
array2[17316]=30'd295074390;
array2[17317]=30'd357913199;
array2[17318]=30'd295074390;
array2[17319]=30'd295074390;
array2[17320]=30'd295074390;
array2[17321]=30'd222764576;
array2[17322]=30'd207191473;
array2[17323]=30'd234504581;
array2[17324]=30'd227165569;
array2[17325]=30'd228216193;
array2[17326]=30'd229266819;
array2[17327]=30'd229266819;
array2[17328]=30'd221916546;
array2[17329]=30'd232392085;
array2[17330]=30'd232392085;
array2[17331]=30'd221916546;
array2[17332]=30'd231362949;
array2[17333]=30'd227159434;
array2[17334]=30'd232392085;
array2[17335]=30'd220861839;
array2[17336]=30'd212454818;
array2[17337]=30'd124307934;
array2[17338]=30'd124307934;
array2[17339]=30'd124307934;
array2[17340]=30'd190356956;
array2[17341]=30'd190356956;
array2[17342]=30'd228181405;
array2[17343]=30'd227159434;
array2[17344]=30'd231362949;
array2[17345]=30'd231362949;
array2[17346]=30'd230317442;
array2[17347]=30'd231362949;
array2[17348]=30'd231364996;
array2[17349]=30'd231362949;
array2[17350]=30'd230317442;
array2[17351]=30'd231364996;
array2[17352]=30'd230317442;
array2[17353]=30'd231362949;
array2[17354]=30'd231362949;
array2[17355]=30'd229266819;
array2[17356]=30'd231362949;
array2[17357]=30'd231362949;
array2[17358]=30'd230317442;
array2[17359]=30'd234504581;
array2[17360]=30'd229266819;
array2[17361]=30'd229266819;
array2[17362]=30'd231362949;
array2[17363]=30'd234504581;
array2[17364]=30'd230317442;
array2[17365]=30'd234504581;
array2[17366]=30'd230317442;
array2[17367]=30'd231362949;
array2[17368]=30'd228212100;
array2[17369]=30'd231364996;
array2[17370]=30'd229266819;
array2[17371]=30'd231362949;
array2[17372]=30'd230317442;
array2[17373]=30'd229266819;
array2[17374]=30'd225072515;
array2[17375]=30'd229266819;
array2[17376]=30'd822672828;
array2[17377]=30'd664345022;
array2[17378]=30'd616102353;
array2[17379]=30'd822672828;
array2[17380]=30'd377085336;
array2[17381]=30'd229270912;
array2[17382]=30'd230317442;
array2[17383]=30'd229270912;
array2[17384]=30'd230317442;
array2[17385]=30'd229266819;
array2[17386]=30'd229266819;
array2[17387]=30'd231362949;
array2[17388]=30'd234504581;
array2[17389]=30'd227165569;
array2[17390]=30'd227165569;
array2[17391]=30'd231362949;
array2[17392]=30'd231362949;
array2[17393]=30'd228216193;
array2[17394]=30'd231362949;
array2[17395]=30'd231362949;
array2[17396]=30'd231362949;
array2[17397]=30'd231359873;
array2[17398]=30'd231362949;
array2[17399]=30'd229266819;
array2[17400]=30'd603537847;
array2[17401]=30'd472496545;
array2[17402]=30'd822672828;
array2[17403]=30'd472496545;
array2[17404]=30'd231362949;
array2[17405]=30'd231362949;
array2[17406]=30'd231362949;
array2[17407]=30'd231362949;
array2[17408]=30'd229266819;
array2[17409]=30'd231362949;
array2[17410]=30'd231362949;
array2[17411]=30'd193577377;
array2[17412]=30'd265736724;
array2[17413]=30'd295074390;
array2[17414]=30'd190356956;
array2[17415]=30'd190356956;
array2[17416]=30'd218607140;
array2[17417]=30'd249001484;
array2[17418]=30'd193577377;
array2[17419]=30'd231362949;
array2[17420]=30'd231364996;
array2[17421]=30'd225072515;
array2[17422]=30'd220861839;
array2[17423]=30'd220861839;
array2[17424]=30'd179916222;
array2[17425]=30'd218607140;
array2[17426]=30'd218607140;
array2[17427]=30'd179916222;
array2[17428]=30'd213516691;
array2[17429]=30'd193577377;
array2[17430]=30'd124307934;
array2[17431]=30'd124307934;
array2[17432]=30'd207191473;
array2[17433]=30'd124307934;
array2[17434]=30'd159912438;
array2[17435]=30'd249001484;
array2[17436]=30'd401997362;
array2[17437]=30'd485780117;
array2[17438]=30'd295074390;
array2[17439]=30'd260631016;
array2[17440]=30'd220861839;
array2[17441]=30'd232392085;
array2[17442]=30'd231362949;
array2[17443]=30'd229266819;
array2[17444]=30'd231364996;
array2[17445]=30'd231362949;
array2[17446]=30'd229266819;
array2[17447]=30'd231362949;
array2[17448]=30'd231362949;
array2[17449]=30'd229266819;
array2[17450]=30'd231364996;
array2[17451]=30'd229266819;
array2[17452]=30'd231362949;
array2[17453]=30'd230317442;
array2[17454]=30'd231362949;
array2[17455]=30'd231362949;
array2[17456]=30'd231362949;
array2[17457]=30'd231362949;
array2[17458]=30'd231362949;
array2[17459]=30'd229266819;
array2[17460]=30'd231362949;
array2[17461]=30'd234504581;
array2[17462]=30'd231362949;
array2[17463]=30'd231362949;
array2[17464]=30'd231362949;
array2[17465]=30'd231362949;
array2[17466]=30'd228216193;
array2[17467]=30'd231362949;
array2[17468]=30'd231362949;
array2[17469]=30'd228216193;
array2[17470]=30'd231362949;
array2[17471]=30'd229266819;
array2[17472]=30'd254365107;
array2[17473]=30'd603537847;
array2[17474]=30'd719920570;
array2[17475]=30'd248105365;
array2[17476]=30'd238691720;
array2[17477]=30'd228216193;
array2[17478]=30'd231364996;
array2[17479]=30'd230317442;
array2[17480]=30'd229266819;
array2[17481]=30'd229266819;
array2[17482]=30'd231362949;
array2[17483]=30'd234504581;
array2[17484]=30'd231359873;
array2[17485]=30'd234499470;
array2[17486]=30'd231362949;
array2[17487]=30'd228216193;
array2[17488]=30'd231362949;
array2[17489]=30'd229266819;
array2[17490]=30'd231362949;
array2[17491]=30'd229266819;
array2[17492]=30'd231359873;
array2[17493]=30'd231364996;
array2[17494]=30'd231362949;
array2[17495]=30'd229266819;
array2[17496]=30'd472496545;
array2[17497]=30'd777593273;
array2[17498]=30'd281654691;
array2[17499]=30'd238691720;
array2[17500]=30'd234504581;
array2[17501]=30'd231359873;
array2[17502]=30'd231362949;
array2[17503]=30'd231362949;
array2[17504]=30'd229266819;
array2[17505]=30'd231362949;
array2[17506]=30'd231362949;
array2[17507]=30'd212454818;
array2[17508]=30'd179916222;
array2[17509]=30'd179916222;
array2[17510]=30'd232392085;
array2[17511]=30'd213516691;
array2[17512]=30'd124307934;
array2[17513]=30'd190356956;
array2[17514]=30'd212454818;
array2[17515]=30'd228181405;
array2[17516]=30'd212454818;
array2[17517]=30'd260631016;
array2[17518]=30'd407216718;
array2[17519]=30'd444954173;
array2[17520]=30'd338018898;
array2[17521]=30'd357913199;
array2[17522]=30'd357913199;
array2[17523]=30'd331763301;
array2[17524]=30'd444954173;
array2[17525]=30'd444954173;
array2[17526]=30'd218607140;
array2[17527]=30'd106464746;
array2[17528]=30'd124307934;
array2[17529]=30'd124307934;
array2[17530]=30'd347490866;
array2[17531]=30'd566515308;
array2[17532]=30'd566515308;
array2[17533]=30'd560184961;
array2[17534]=30'd560184961;
array2[17535]=30'd485780117;
array2[17536]=30'd331763301;
array2[17537]=30'd260631016;
array2[17538]=30'd212454818;
array2[17539]=30'd221916546;
array2[17540]=30'd228216193;
array2[17541]=30'd230317442;
array2[17542]=30'd230317442;
array2[17543]=30'd229266819;
array2[17544]=30'd228216193;
array2[17545]=30'd228216193;
array2[17546]=30'd230317442;
array2[17547]=30'd230317442;
array2[17548]=30'd229270912;
array2[17549]=30'd229266819;
array2[17550]=30'd231362949;
array2[17551]=30'd230317442;
array2[17552]=30'd231362949;
array2[17553]=30'd234504581;
array2[17554]=30'd231362949;
array2[17555]=30'd231364996;
array2[17556]=30'd234504581;
array2[17557]=30'd229266819;
array2[17558]=30'd230317442;
array2[17559]=30'd231362949;
array2[17560]=30'd234504581;
array2[17561]=30'd229266819;
array2[17562]=30'd231362949;
array2[17563]=30'd229270912;
array2[17564]=30'd227165569;
array2[17565]=30'd227159434;
array2[17566]=30'd230317442;
array2[17567]=30'd230317442;
array2[17568]=30'd212454818;
array2[17569]=30'd256519562;
array2[17570]=30'd256519562;
array2[17571]=30'd234504581;
array2[17572]=30'd228216193;
array2[17573]=30'd228216193;
array2[17574]=30'd228212100;
array2[17575]=30'd229266819;
array2[17576]=30'd231362949;
array2[17577]=30'd231359873;
array2[17578]=30'd229266819;
array2[17579]=30'd229266819;
array2[17580]=30'd231362949;
array2[17581]=30'd229270912;
array2[17582]=30'd231364996;
array2[17583]=30'd231362949;
array2[17584]=30'd231359873;
array2[17585]=30'd228216193;
array2[17586]=30'd231364996;
array2[17587]=30'd231364996;
array2[17588]=30'd232417668;
array2[17589]=30'd230317442;
array2[17590]=30'd231364996;
array2[17591]=30'd230317442;
array2[17592]=30'd256519562;
array2[17593]=30'd256519562;
array2[17594]=30'd234499470;
array2[17595]=30'd234504581;
array2[17596]=30'd228212100;
array2[17597]=30'd234504581;
array2[17598]=30'd234504581;
array2[17599]=30'd231362949;
array2[17600]=30'd231364996;
array2[17601]=30'd229266819;
array2[17602]=30'd229266819;
array2[17603]=30'd231362949;
array2[17604]=30'd231359873;
array2[17605]=30'd234504581;
array2[17606]=30'd231362949;
array2[17607]=30'd195647926;
array2[17608]=30'd299264555;
array2[17609]=30'd331763301;
array2[17610]=30'd299264555;
array2[17611]=30'd265736724;
array2[17612]=30'd483727963;
array2[17613]=30'd645112409;
array2[17614]=30'd819020415;
array2[17615]=30'd828452495;
array2[17616]=30'd560184961;
array2[17617]=30'd375721588;
array2[17618]=30'd375721588;
array2[17619]=30'd518272648;
array2[17620]=30'd819020415;
array2[17621]=30'd819020415;
array2[17622]=30'd606320275;
array2[17623]=30'd249001484;
array2[17624]=30'd106464746;
array2[17625]=30'd83428824;
array2[17626]=30'd449120871;
array2[17627]=30'd770812573;
array2[17628]=30'd799112870;
array2[17629]=30'd678602388;
array2[17630]=30'd606320275;
array2[17631]=30'd518272648;
array2[17632]=30'd560184961;
array2[17633]=30'd481587821;
array2[17634]=30'd375721588;
array2[17635]=30'd260631016;
array2[17636]=30'd231362949;
array2[17637]=30'd231362949;
array2[17638]=30'd231364996;
array2[17639]=30'd231362949;
array2[17640]=30'd229266819;
array2[17641]=30'd231362949;
array2[17642]=30'd231362949;
array2[17643]=30'd229266819;
array2[17644]=30'd231362949;
array2[17645]=30'd231362949;
array2[17646]=30'd231362949;
array2[17647]=30'd230317442;
array2[17648]=30'd231364996;
array2[17649]=30'd228216193;
array2[17650]=30'd231362949;
array2[17651]=30'd231362949;
array2[17652]=30'd231362949;
array2[17653]=30'd229266819;
array2[17654]=30'd229266819;
array2[17655]=30'd231362949;
array2[17656]=30'd229266819;
array2[17657]=30'd230317442;
array2[17658]=30'd231362949;
array2[17659]=30'd231362949;
array2[17660]=30'd228216193;
array2[17661]=30'd230317442;
array2[17662]=30'd229270912;
array2[17663]=30'd229266819;
array2[17664]=30'd212454818;
array2[17665]=30'd231359873;
array2[17666]=30'd227165569;
array2[17667]=30'd234504581;
array2[17668]=30'd240774546;
array2[17669]=30'd232392085;
array2[17670]=30'd232392085;
array2[17671]=30'd232392085;
array2[17672]=30'd232392085;
array2[17673]=30'd232392085;
array2[17674]=30'd232392085;
array2[17675]=30'd234499470;
array2[17676]=30'd234499470;
array2[17677]=30'd236604812;
array2[17678]=30'd232392085;
array2[17679]=30'd234504581;
array2[17680]=30'd229270912;
array2[17681]=30'd231364996;
array2[17682]=30'd229270912;
array2[17683]=30'd232422779;
array2[17684]=30'd229270912;
array2[17685]=30'd231364996;
array2[17686]=30'd229270912;
array2[17687]=30'd231364996;
array2[17688]=30'd231362949;
array2[17689]=30'd231362949;
array2[17690]=30'd228216193;
array2[17691]=30'd238691720;
array2[17692]=30'd232392085;
array2[17693]=30'd232392085;
array2[17694]=30'd232392085;
array2[17695]=30'd227159434;
array2[17696]=30'd232392085;
array2[17697]=30'd227159434;
array2[17698]=30'd234499470;
array2[17699]=30'd234499470;
array2[17700]=30'd234499470;
array2[17701]=30'd232392085;
array2[17702]=30'd232392085;
array2[17703]=30'd124307934;
array2[17704]=30'd218607140;
array2[17705]=30'd265736724;
array2[17706]=30'd295074390;
array2[17707]=30'd560184961;
array2[17708]=30'd768729747;
array2[17709]=30'd851505800;
array2[17710]=30'd865130113;
array2[17711]=30'd865130113;
array2[17712]=30'd606320275;
array2[17713]=30'd375721588;
array2[17714]=30'd375721588;
array2[17715]=30'd566515308;
array2[17716]=30'd851505800;
array2[17717]=30'd858839683;
array2[17718]=30'd828452495;
array2[17719]=30'd407216718;
array2[17720]=30'd159912438;
array2[17721]=30'd106464746;
array2[17722]=30'd319215128;
array2[17723]=30'd672348794;
array2[17724]=30'd858839683;
array2[17725]=30'd828452495;
array2[17726]=30'd799112870;
array2[17727]=30'd678602388;
array2[17728]=30'd606320275;
array2[17729]=30'd518272648;
array2[17730]=30'd539218630;
array2[17731]=30'd450208341;
array2[17732]=30'd179916222;
array2[17733]=30'd195647926;
array2[17734]=30'd227159434;
array2[17735]=30'd228216193;
array2[17736]=30'd228216193;
array2[17737]=30'd230317442;
array2[17738]=30'd231362949;
array2[17739]=30'd231364996;
array2[17740]=30'd231362949;
array2[17741]=30'd229266819;
array2[17742]=30'd231362949;
array2[17743]=30'd230317442;
array2[17744]=30'd231362949;
array2[17745]=30'd229266819;
array2[17746]=30'd231362949;
array2[17747]=30'd231362949;
array2[17748]=30'd229266819;
array2[17749]=30'd231362949;
array2[17750]=30'd231362949;
array2[17751]=30'd231362949;
array2[17752]=30'd231362949;
array2[17753]=30'd231362949;
array2[17754]=30'd229266819;
array2[17755]=30'd231362949;
array2[17756]=30'd231362949;
array2[17757]=30'd231364996;
array2[17758]=30'd231362949;
array2[17759]=30'd231362949;
array2[17760]=30'd260631016;
array2[17761]=30'd280568333;
array2[17762]=30'd280568333;
array2[17763]=30'd307771998;
array2[17764]=30'd390446940;
array2[17765]=30'd461700935;
array2[17766]=30'd461700935;
array2[17767]=30'd461700935;
array2[17768]=30'd461700935;
array2[17769]=30'd461700935;
array2[17770]=30'd461700935;
array2[17771]=30'd461700935;
array2[17772]=30'd461700935;
array2[17773]=30'd461700935;
array2[17774]=30'd461700935;
array2[17775]=30'd328674981;
array2[17776]=30'd280568333;
array2[17777]=30'd280568333;
array2[17778]=30'd280568333;
array2[17779]=30'd280568333;
array2[17780]=30'd280568333;
array2[17781]=30'd280568333;
array2[17782]=30'd280568333;
array2[17783]=30'd280568333;
array2[17784]=30'd280568333;
array2[17785]=30'd280568333;
array2[17786]=30'd280568333;
array2[17787]=30'd395649781;
array2[17788]=30'd461700935;
array2[17789]=30'd461700935;
array2[17790]=30'd461700935;
array2[17791]=30'd461700935;
array2[17792]=30'd461700935;
array2[17793]=30'd461700935;
array2[17794]=30'd461700935;
array2[17795]=30'd461700935;
array2[17796]=30'd461700935;
array2[17797]=30'd461700935;
array2[17798]=30'd357996288;
array2[17799]=30'd218607140;
array2[17800]=30'd218607140;
array2[17801]=30'd218607140;
array2[17802]=30'd434416250;
array2[17803]=30'd768729747;
array2[17804]=30'd828452495;
array2[17805]=30'd851505800;
array2[17806]=30'd858839683;
array2[17807]=30'd858839683;
array2[17808]=30'd606320275;
array2[17809]=30'd375721588;
array2[17810]=30'd375721588;
array2[17811]=30'd560184961;
array2[17812]=30'd851505800;
array2[17813]=30'd851505800;
array2[17814]=30'd851505800;
array2[17815]=30'd506770009;
array2[17816]=30'd295074390;
array2[17817]=30'd131612152;
array2[17818]=30'd106464746;
array2[17819]=30'd566515308;
array2[17820]=30'd828452495;
array2[17821]=30'd851505800;
array2[17822]=30'd851505800;
array2[17823]=30'd851505800;
array2[17824]=30'd768729747;
array2[17825]=30'd678602388;
array2[17826]=30'd560184961;
array2[17827]=30'd481587821;
array2[17828]=30'd401997362;
array2[17829]=30'd383147560;
array2[17830]=30'd179916222;
array2[17831]=30'd179916222;
array2[17832]=30'd212454818;
array2[17833]=30'd228212100;
array2[17834]=30'd231362949;
array2[17835]=30'd231362949;
array2[17836]=30'd231362949;
array2[17837]=30'd229266819;
array2[17838]=30'd231362949;
array2[17839]=30'd231362949;
array2[17840]=30'd231364996;
array2[17841]=30'd230317442;
array2[17842]=30'd231362949;
array2[17843]=30'd229266819;
array2[17844]=30'd228216193;
array2[17845]=30'd231364996;
array2[17846]=30'd231364996;
array2[17847]=30'd231362949;
array2[17848]=30'd231362949;
array2[17849]=30'd231362949;
array2[17850]=30'd231362949;
array2[17851]=30'd231362949;
array2[17852]=30'd231362949;
array2[17853]=30'd229266819;
array2[17854]=30'd234504581;
array2[17855]=30'd230317442;
array2[17856]=30'd390446940;
array2[17857]=30'd409311115;
array2[17858]=30'd409311115;
array2[17859]=30'd409311115;
array2[17860]=30'd429185963;
array2[17861]=30'd423950257;
array2[17862]=30'd426044336;
array2[17863]=30'd423950257;
array2[17864]=30'd426044336;
array2[17865]=30'd423950257;
array2[17866]=30'd423950257;
array2[17867]=30'd426044336;
array2[17868]=30'd423950257;
array2[17869]=30'd426044336;
array2[17870]=30'd426044336;
array2[17871]=30'd429185963;
array2[17872]=30'd409311115;
array2[17873]=30'd409311115;
array2[17874]=30'd409311115;
array2[17875]=30'd409311115;
array2[17876]=30'd409311115;
array2[17877]=30'd409311115;
array2[17878]=30'd409311115;
array2[17879]=30'd409311115;
array2[17880]=30'd409311115;
array2[17881]=30'd409311115;
array2[17882]=30'd409311115;
array2[17883]=30'd429185963;
array2[17884]=30'd426044336;
array2[17885]=30'd426044336;
array2[17886]=30'd423950257;
array2[17887]=30'd426044336;
array2[17888]=30'd426044336;
array2[17889]=30'd426044336;
array2[17890]=30'd423950257;
array2[17891]=30'd426044336;
array2[17892]=30'd423950257;
array2[17893]=30'd426044336;
array2[17894]=30'd429185963;
array2[17895]=30'd409311115;
array2[17896]=30'd395649781;
array2[17897]=30'd434416250;
array2[17898]=30'd770812573;
array2[17899]=30'd851505800;
array2[17900]=30'd851505800;
array2[17901]=30'd858839683;
array2[17902]=30'd865130113;
array2[17903]=30'd865130113;
array2[17904]=30'd606320275;
array2[17905]=30'd375721588;
array2[17906]=30'd434416250;
array2[17907]=30'd713179821;
array2[17908]=30'd858839683;
array2[17909]=30'd851505800;
array2[17910]=30'd851505800;
array2[17911]=30'd518272648;
array2[17912]=30'd375721588;
array2[17913]=30'd295074390;
array2[17914]=30'd159912438;
array2[17915]=30'd518272648;
array2[17916]=30'd770816666;
array2[17917]=30'd770816666;
array2[17918]=30'd799112870;
array2[17919]=30'd851505800;
array2[17920]=30'd851505800;
array2[17921]=30'd828452495;
array2[17922]=30'd770812573;
array2[17923]=30'd518272648;
array2[17924]=30'd481587821;
array2[17925]=30'd711090860;
array2[17926]=30'd768729747;
array2[17927]=30'd727851632;
array2[17928]=30'd401997362;
array2[17929]=30'd190356956;
array2[17930]=30'd213516691;
array2[17931]=30'd230307208;
array2[17932]=30'd231364996;
array2[17933]=30'd229270912;
array2[17934]=30'd229266819;
array2[17935]=30'd229266819;
array2[17936]=30'd231362949;
array2[17937]=30'd231362949;
array2[17938]=30'd234504581;
array2[17939]=30'd227165569;
array2[17940]=30'd234504581;
array2[17941]=30'd231362949;
array2[17942]=30'd231362949;
array2[17943]=30'd231362949;
array2[17944]=30'd231362949;
array2[17945]=30'd229266819;
array2[17946]=30'd231359873;
array2[17947]=30'd231362949;
array2[17948]=30'd231362949;
array2[17949]=30'd229266819;
array2[17950]=30'd230317442;
array2[17951]=30'd229270912;
array2[17952]=30'd409311115;
array2[17953]=30'd426044336;
array2[17954]=30'd426044336;
array2[17955]=30'd426044336;
array2[17956]=30'd426044336;
array2[17957]=30'd426044336;
array2[17958]=30'd426044336;
array2[17959]=30'd426044336;
array2[17960]=30'd426044336;
array2[17961]=30'd426044336;
array2[17962]=30'd426044336;
array2[17963]=30'd426044336;
array2[17964]=30'd423950257;
array2[17965]=30'd423950257;
array2[17966]=30'd426044336;
array2[17967]=30'd426044336;
array2[17968]=30'd426044336;
array2[17969]=30'd426044336;
array2[17970]=30'd423950257;
array2[17971]=30'd423950257;
array2[17972]=30'd423950257;
array2[17973]=30'd423950257;
array2[17974]=30'd423950257;
array2[17975]=30'd426044336;
array2[17976]=30'd423950257;
array2[17977]=30'd423950257;
array2[17978]=30'd426044336;
array2[17979]=30'd423950257;
array2[17980]=30'd426044336;
array2[17981]=30'd426044336;
array2[17982]=30'd426044336;
array2[17983]=30'd426044336;
array2[17984]=30'd426044336;
array2[17985]=30'd426044336;
array2[17986]=30'd426044336;
array2[17987]=30'd426044336;
array2[17988]=30'd426044336;
array2[17989]=30'd423950257;
array2[17990]=30'd423950257;
array2[17991]=30'd461700935;
array2[17992]=30'd375721588;
array2[17993]=30'd770816666;
array2[17994]=30'd851505800;
array2[17995]=30'd851505800;
array2[17996]=30'd858839683;
array2[17997]=30'd865130113;
array2[17998]=30'd858839683;
array2[17999]=30'd851505800;
array2[18000]=30'd631447172;
array2[18001]=30'd375721588;
array2[18002]=30'd434416250;
array2[18003]=30'd819020415;
array2[18004]=30'd851505800;
array2[18005]=30'd851505800;
array2[18006]=30'd851505800;
array2[18007]=30'd518272648;
array2[18008]=30'd375721588;
array2[18009]=30'd357913199;
array2[18010]=30'd566515308;
array2[18011]=30'd631447172;
array2[18012]=30'd631447172;
array2[18013]=30'd713179821;
array2[18014]=30'd732038833;
array2[18015]=30'd819020415;
array2[18016]=30'd851505800;
array2[18017]=30'd858839683;
array2[18018]=30'd851505800;
array2[18019]=30'd828452495;
array2[18020]=30'd770812573;
array2[18021]=30'd678602388;
array2[18022]=30'd851505800;
array2[18023]=30'd851505800;
array2[18024]=30'd819020415;
array2[18025]=30'd713179821;
array2[18026]=30'd347490866;
array2[18027]=30'd190356956;
array2[18028]=30'd221916546;
array2[18029]=30'd231362949;
array2[18030]=30'd230317442;
array2[18031]=30'd231362949;
array2[18032]=30'd231364996;
array2[18033]=30'd231362949;
array2[18034]=30'd231362949;
array2[18035]=30'd231362949;
array2[18036]=30'd231362949;
array2[18037]=30'd231362949;
array2[18038]=30'd231362949;
array2[18039]=30'd234504581;
array2[18040]=30'd231362949;
array2[18041]=30'd231362949;
array2[18042]=30'd230317442;
array2[18043]=30'd229266819;
array2[18044]=30'd231362949;
array2[18045]=30'd231362949;
array2[18046]=30'd231362949;
array2[18047]=30'd231362949;
array2[18048]=30'd409311115;
array2[18049]=30'd426044336;
array2[18050]=30'd426044336;
array2[18051]=30'd493111164;
array2[18052]=30'd635645720;
array2[18053]=30'd672324351;
array2[18054]=30'd672324351;
array2[18055]=30'd672324351;
array2[18056]=30'd672324351;
array2[18057]=30'd672324351;
array2[18058]=30'd672324351;
array2[18059]=30'd672324351;
array2[18060]=30'd672324351;
array2[18061]=30'd672324351;
array2[18062]=30'd672324351;
array2[18063]=30'd493111164;
array2[18064]=30'd426044336;
array2[18065]=30'd435467177;
array2[18066]=30'd426044336;
array2[18067]=30'd426044336;
array2[18068]=30'd426044336;
array2[18069]=30'd426044336;
array2[18070]=30'd426044336;
array2[18071]=30'd426044336;
array2[18072]=30'd426044336;
array2[18073]=30'd426044336;
array2[18074]=30'd435467177;
array2[18075]=30'd582196031;
array2[18076]=30'd672324351;
array2[18077]=30'd672324351;
array2[18078]=30'd672324351;
array2[18079]=30'd672324351;
array2[18080]=30'd672324351;
array2[18081]=30'd672324351;
array2[18082]=30'd672324351;
array2[18083]=30'd718417640;
array2[18084]=30'd672324351;
array2[18085]=30'd672324351;
array2[18086]=30'd582196031;
array2[18087]=30'd395649781;
array2[18088]=30'd566515308;
array2[18089]=30'd851505800;
array2[18090]=30'd851505800;
array2[18091]=30'd851505800;
array2[18092]=30'd851505800;
array2[18093]=30'd858839683;
array2[18094]=30'd858839683;
array2[18095]=30'd851505800;
array2[18096]=30'd828452495;
array2[18097]=30'd631447172;
array2[18098]=30'd565444213;
array2[18099]=30'd828452495;
array2[18100]=30'd865130113;
array2[18101]=30'd865130113;
array2[18102]=30'd858839683;
array2[18103]=30'd606320275;
array2[18104]=30'd375721588;
array2[18105]=30'd375721588;
array2[18106]=30'd631447172;
array2[18107]=30'd799112870;
array2[18108]=30'd672348794;
array2[18109]=30'd566515308;
array2[18110]=30'd672348794;
array2[18111]=30'd711090860;
array2[18112]=30'd770812573;
array2[18113]=30'd828452495;
array2[18114]=30'd858839683;
array2[18115]=30'd858839683;
array2[18116]=30'd865130113;
array2[18117]=30'd858839683;
array2[18118]=30'd858839683;
array2[18119]=30'd865130113;
array2[18120]=30'd858839683;
array2[18121]=30'd858839683;
array2[18122]=30'd828452495;
array2[18123]=30'd677571193;
array2[18124]=30'd179916222;
array2[18125]=30'd231364996;
array2[18126]=30'd228216193;
array2[18127]=30'd231362949;
array2[18128]=30'd231364996;
array2[18129]=30'd229266819;
array2[18130]=30'd229266819;
array2[18131]=30'd231362949;
array2[18132]=30'd231362949;
array2[18133]=30'd234504581;
array2[18134]=30'd234504581;
array2[18135]=30'd234504581;
array2[18136]=30'd231359873;
array2[18137]=30'd231362949;
array2[18138]=30'd229266819;
array2[18139]=30'd229266819;
array2[18140]=30'd230317442;
array2[18141]=30'd229266819;
array2[18142]=30'd234504581;
array2[18143]=30'd231364996;
array2[18144]=30'd646169309;
array2[18145]=30'd672324351;
array2[18146]=30'd672324351;
array2[18147]=30'd672324351;
array2[18148]=30'd718417640;
array2[18149]=30'd728897252;
array2[18150]=30'd728897252;
array2[18151]=30'd728897252;
array2[18152]=30'd728897252;
array2[18153]=30'd728897252;
array2[18154]=30'd728897252;
array2[18155]=30'd728897252;
array2[18156]=30'd728897252;
array2[18157]=30'd728897252;
array2[18158]=30'd728897252;
array2[18159]=30'd718417640;
array2[18160]=30'd672324351;
array2[18161]=30'd718417640;
array2[18162]=30'd718417640;
array2[18163]=30'd718417640;
array2[18164]=30'd718417640;
array2[18165]=30'd718417640;
array2[18166]=30'd672324351;
array2[18167]=30'd718417640;
array2[18168]=30'd672324351;
array2[18169]=30'd672324351;
array2[18170]=30'd672324351;
array2[18171]=30'd718417640;
array2[18172]=30'd728897252;
array2[18173]=30'd728897252;
array2[18174]=30'd728897252;
array2[18175]=30'd728897252;
array2[18176]=30'd728897252;
array2[18177]=30'd728897252;
array2[18178]=30'd728897252;
array2[18179]=30'd728897252;
array2[18180]=30'd728897252;
array2[18181]=30'd728897252;
array2[18182]=30'd646169309;
array2[18183]=30'd299264555;
array2[18184]=30'd799112870;
array2[18185]=30'd858839683;
array2[18186]=30'd851505800;
array2[18187]=30'd858839683;
array2[18188]=30'd858839683;
array2[18189]=30'd865130113;
array2[18190]=30'd865130113;
array2[18191]=30'd865130113;
array2[18192]=30'd858839683;
array2[18193]=30'd865130113;
array2[18194]=30'd865130113;
array2[18195]=30'd865130113;
array2[18196]=30'd865130113;
array2[18197]=30'd858839683;
array2[18198]=30'd858839683;
array2[18199]=30'd672348794;
array2[18200]=30'd434416250;
array2[18201]=30'd481587821;
array2[18202]=30'd711090860;
array2[18203]=30'd865130113;
array2[18204]=30'd828452495;
array2[18205]=30'd711090860;
array2[18206]=30'd606320275;
array2[18207]=30'd604201637;
array2[18208]=30'd711090860;
array2[18209]=30'd768729747;
array2[18210]=30'd828452495;
array2[18211]=30'd858839683;
array2[18212]=30'd865130113;
array2[18213]=30'd851505800;
array2[18214]=30'd865130113;
array2[18215]=30'd858839683;
array2[18216]=30'd858839683;
array2[18217]=30'd858839683;
array2[18218]=30'd858839683;
array2[18219]=30'd764529268;
array2[18220]=30'd383147560;
array2[18221]=30'd213516691;
array2[18222]=30'd231362949;
array2[18223]=30'd229266819;
array2[18224]=30'd228216193;
array2[18225]=30'd229266819;
array2[18226]=30'd231364996;
array2[18227]=30'd229266819;
array2[18228]=30'd231364996;
array2[18229]=30'd231362949;
array2[18230]=30'd230317442;
array2[18231]=30'd231362949;
array2[18232]=30'd229266819;
array2[18233]=30'd231362949;
array2[18234]=30'd231362949;
array2[18235]=30'd231362949;
array2[18236]=30'd231362949;
array2[18237]=30'd229266819;
array2[18238]=30'd231362949;
array2[18239]=30'd227165569;
array2[18240]=30'd713202349;
array2[18241]=30'd728897252;
array2[18242]=30'd728897252;
array2[18243]=30'd728897252;
array2[18244]=30'd728897252;
array2[18245]=30'd728897252;
array2[18246]=30'd728897252;
array2[18247]=30'd728897252;
array2[18248]=30'd728897252;
array2[18249]=30'd728897252;
array2[18250]=30'd728897252;
array2[18251]=30'd728897252;
array2[18252]=30'd728897252;
array2[18253]=30'd728897252;
array2[18254]=30'd728897252;
array2[18255]=30'd728897252;
array2[18256]=30'd728897252;
array2[18257]=30'd728897252;
array2[18258]=30'd728897252;
array2[18259]=30'd728897252;
array2[18260]=30'd728897252;
array2[18261]=30'd728897252;
array2[18262]=30'd728897252;
array2[18263]=30'd728897252;
array2[18264]=30'd728897252;
array2[18265]=30'd728897252;
array2[18266]=30'd728897252;
array2[18267]=30'd728897252;
array2[18268]=30'd728897252;
array2[18269]=30'd728897252;
array2[18270]=30'd728897252;
array2[18271]=30'd728897252;
array2[18272]=30'd728897252;
array2[18273]=30'd728897252;
array2[18274]=30'd728897252;
array2[18275]=30'd728897252;
array2[18276]=30'd728897252;
array2[18277]=30'd718417640;
array2[18278]=30'd481587821;
array2[18279]=30'd606320275;
array2[18280]=30'd851505800;
array2[18281]=30'd858839683;
array2[18282]=30'd865130113;
array2[18283]=30'd851505800;
array2[18284]=30'd865130113;
array2[18285]=30'd865130113;
array2[18286]=30'd858839683;
array2[18287]=30'd858839683;
array2[18288]=30'd858839683;
array2[18289]=30'd858839683;
array2[18290]=30'd858839683;
array2[18291]=30'd858839683;
array2[18292]=30'd858839683;
array2[18293]=30'd858839683;
array2[18294]=30'd858839683;
array2[18295]=30'd828452495;
array2[18296]=30'd727851632;
array2[18297]=30'd764529268;
array2[18298]=30'd851505800;
array2[18299]=30'd865130113;
array2[18300]=30'd865130113;
array2[18301]=30'd858839683;
array2[18302]=30'd828452495;
array2[18303]=30'd828452495;
array2[18304]=30'd768729747;
array2[18305]=30'd819020415;
array2[18306]=30'd851505800;
array2[18307]=30'd865130113;
array2[18308]=30'd858839683;
array2[18309]=30'd865130113;
array2[18310]=30'd865130113;
array2[18311]=30'd858839683;
array2[18312]=30'd858839683;
array2[18313]=30'd858839683;
array2[18314]=30'd858839683;
array2[18315]=30'd851505800;
array2[18316]=30'd713179821;
array2[18317]=30'd401997362;
array2[18318]=30'd212454818;
array2[18319]=30'd234504581;
array2[18320]=30'd228212100;
array2[18321]=30'd229266819;
array2[18322]=30'd231362949;
array2[18323]=30'd231362949;
array2[18324]=30'd231364996;
array2[18325]=30'd231362949;
array2[18326]=30'd231359873;
array2[18327]=30'd227165569;
array2[18328]=30'd231362949;
array2[18329]=30'd229266819;
array2[18330]=30'd231362949;
array2[18331]=30'd228216193;
array2[18332]=30'd228216193;
array2[18333]=30'd231359873;
array2[18334]=30'd231362949;
array2[18335]=30'd231362949;
array2[18336]=30'd711090860;
array2[18337]=30'd728897252;
array2[18338]=30'd728897252;
array2[18339]=30'd758240964;
array2[18340]=30'd828452495;
array2[18341]=30'd865130113;
array2[18342]=30'd865130113;
array2[18343]=30'd865130113;
array2[18344]=30'd865130113;
array2[18345]=30'd865130113;
array2[18346]=30'd865130113;
array2[18347]=30'd865130113;
array2[18348]=30'd865130113;
array2[18349]=30'd865130113;
array2[18350]=30'd865130113;
array2[18351]=30'd758240964;
array2[18352]=30'd728897252;
array2[18353]=30'd728897252;
array2[18354]=30'd728897252;
array2[18355]=30'd728897252;
array2[18356]=30'd728897252;
array2[18357]=30'd728897252;
array2[18358]=30'd728897252;
array2[18359]=30'd728897252;
array2[18360]=30'd728897252;
array2[18361]=30'd728897252;
array2[18362]=30'd728897252;
array2[18363]=30'd828452495;
array2[18364]=30'd865130113;
array2[18365]=30'd865130113;
array2[18366]=30'd865130113;
array2[18367]=30'd865130113;
array2[18368]=30'd865130113;
array2[18369]=30'd865130113;
array2[18370]=30'd865130113;
array2[18371]=30'd865130113;
array2[18372]=30'd865130113;
array2[18373]=30'd819020415;
array2[18374]=30'd347490866;
array2[18375]=30'd770816666;
array2[18376]=30'd851505800;
array2[18377]=30'd851505800;
array2[18378]=30'd858839683;
array2[18379]=30'd858839683;
array2[18380]=30'd865130113;
array2[18381]=30'd865130113;
array2[18382]=30'd858839683;
array2[18383]=30'd858839683;
array2[18384]=30'd865130113;
array2[18385]=30'd865130113;
array2[18386]=30'd858839683;
array2[18387]=30'd858839683;
array2[18388]=30'd858839683;
array2[18389]=30'd858839683;
array2[18390]=30'd858839683;
array2[18391]=30'd858839683;
array2[18392]=30'd858839683;
array2[18393]=30'd858839683;
array2[18394]=30'd858839683;
array2[18395]=30'd858839683;
array2[18396]=30'd858839683;
array2[18397]=30'd858839683;
array2[18398]=30'd858839683;
array2[18399]=30'd858839683;
array2[18400]=30'd858839683;
array2[18401]=30'd858839683;
array2[18402]=30'd858839683;
array2[18403]=30'd858839683;
array2[18404]=30'd858839683;
array2[18405]=30'd858839683;
array2[18406]=30'd858839683;
array2[18407]=30'd865130113;
array2[18408]=30'd858839683;
array2[18409]=30'd858839683;
array2[18410]=30'd828452495;
array2[18411]=30'd828452495;
array2[18412]=30'd828452495;
array2[18413]=30'd506770009;
array2[18414]=30'd207191473;
array2[18415]=30'd234504581;
array2[18416]=30'd228212100;
array2[18417]=30'd231359873;
array2[18418]=30'd231362949;
array2[18419]=30'd231362949;
array2[18420]=30'd231362949;
array2[18421]=30'd228216193;
array2[18422]=30'd231359873;
array2[18423]=30'd231362949;
array2[18424]=30'd231362949;
array2[18425]=30'd231362949;
array2[18426]=30'd234504581;
array2[18427]=30'd227165569;
array2[18428]=30'd231362949;
array2[18429]=30'd231362949;
array2[18430]=30'd231362949;
array2[18431]=30'd229266819;
array2[18432]=30'd823228019;
array2[18433]=30'd865130113;
array2[18434]=30'd865130113;
array2[18435]=30'd865130113;
array2[18436]=30'd906004072;
array2[18437]=30'd906004072;
array2[18438]=30'd906004072;
array2[18439]=30'd906004072;
array2[18440]=30'd906004072;
array2[18441]=30'd906004072;
array2[18442]=30'd906004072;
array2[18443]=30'd906004072;
array2[18444]=30'd906004072;
array2[18445]=30'd906004072;
array2[18446]=30'd906004072;
array2[18447]=30'd865130113;
array2[18448]=30'd865130113;
array2[18449]=30'd865130113;
array2[18450]=30'd865130113;
array2[18451]=30'd865130113;
array2[18452]=30'd865130113;
array2[18453]=30'd865130113;
array2[18454]=30'd865130113;
array2[18455]=30'd865130113;
array2[18456]=30'd865130113;
array2[18457]=30'd865130113;
array2[18458]=30'd865130113;
array2[18459]=30'd906004072;
array2[18460]=30'd906004072;
array2[18461]=30'd906004072;
array2[18462]=30'd906004072;
array2[18463]=30'd906004072;
array2[18464]=30'd906004072;
array2[18465]=30'd906004072;
array2[18466]=30'd906004072;
array2[18467]=30'd906004072;
array2[18468]=30'd906004072;
array2[18469]=30'd865130113;
array2[18470]=30'd347490866;
array2[18471]=30'd819020415;
array2[18472]=30'd858839683;
array2[18473]=30'd858839683;
array2[18474]=30'd858839683;
array2[18475]=30'd851505800;
array2[18476]=30'd858839683;
array2[18477]=30'd858839683;
array2[18478]=30'd858839683;
array2[18479]=30'd858839683;
array2[18480]=30'd858839683;
array2[18481]=30'd858839683;
array2[18482]=30'd858839683;
array2[18483]=30'd858839683;
array2[18484]=30'd858839683;
array2[18485]=30'd858839683;
array2[18486]=30'd858839683;
array2[18487]=30'd858839683;
array2[18488]=30'd858839683;
array2[18489]=30'd858839683;
array2[18490]=30'd858839683;
array2[18491]=30'd858839683;
array2[18492]=30'd858839683;
array2[18493]=30'd858839683;
array2[18494]=30'd858839683;
array2[18495]=30'd858839683;
array2[18496]=30'd865130113;
array2[18497]=30'd865130113;
array2[18498]=30'd858839683;
array2[18499]=30'd858839683;
array2[18500]=30'd858839683;
array2[18501]=30'd858839683;
array2[18502]=30'd865130113;
array2[18503]=30'd865130113;
array2[18504]=30'd858839683;
array2[18505]=30'd819020415;
array2[18506]=30'd444954173;
array2[18507]=30'd538207812;
array2[18508]=30'd851505800;
array2[18509]=30'd538207812;
array2[18510]=30'd186252693;
array2[18511]=30'd229270912;
array2[18512]=30'd231362949;
array2[18513]=30'd229270912;
array2[18514]=30'd232417668;
array2[18515]=30'd231362949;
array2[18516]=30'd231362949;
array2[18517]=30'd231362949;
array2[18518]=30'd231359873;
array2[18519]=30'd231359873;
array2[18520]=30'd231362949;
array2[18521]=30'd231362949;
array2[18522]=30'd234504581;
array2[18523]=30'd228216193;
array2[18524]=30'd228216193;
array2[18525]=30'd231362949;
array2[18526]=30'd231362949;
array2[18527]=30'd231362949;
array2[18528]=30'd823228019;
array2[18529]=30'd906004072;
array2[18530]=30'd906004072;
array2[18531]=30'd906004072;
array2[18532]=30'd906004072;
array2[18533]=30'd906004072;
array2[18534]=30'd906004072;
array2[18535]=30'd906004072;
array2[18536]=30'd906004072;
array2[18537]=30'd906004072;
array2[18538]=30'd906004072;
array2[18539]=30'd906004072;
array2[18540]=30'd906004072;
array2[18541]=30'd906004072;
array2[18542]=30'd906004072;
array2[18543]=30'd906004072;
array2[18544]=30'd906004072;
array2[18545]=30'd906004072;
array2[18546]=30'd906004072;
array2[18547]=30'd906004072;
array2[18548]=30'd906004072;
array2[18549]=30'd906004072;
array2[18550]=30'd906004072;
array2[18551]=30'd906004072;
array2[18552]=30'd906004072;
array2[18553]=30'd906004072;
array2[18554]=30'd906004072;
array2[18555]=30'd906004072;
array2[18556]=30'd906004072;
array2[18557]=30'd906004072;
array2[18558]=30'd906004072;
array2[18559]=30'd906004072;
array2[18560]=30'd906004072;
array2[18561]=30'd906004072;
array2[18562]=30'd906004072;
array2[18563]=30'd906004072;
array2[18564]=30'd906004072;
array2[18565]=30'd823228019;
array2[18566]=30'd352736774;
array2[18567]=30'd819020415;
array2[18568]=30'd858839683;
array2[18569]=30'd865130113;
array2[18570]=30'd858839683;
array2[18571]=30'd858839683;
array2[18572]=30'd865130113;
array2[18573]=30'd858839683;
array2[18574]=30'd858839683;
array2[18575]=30'd858839683;
array2[18576]=30'd858839683;
array2[18577]=30'd858839683;
array2[18578]=30'd858839683;
array2[18579]=30'd858839683;
array2[18580]=30'd858839683;
array2[18581]=30'd858839683;
array2[18582]=30'd858839683;
array2[18583]=30'd865130113;
array2[18584]=30'd865130113;
array2[18585]=30'd858839683;
array2[18586]=30'd858839683;
array2[18587]=30'd858839683;
array2[18588]=30'd858839683;
array2[18589]=30'd858839683;
array2[18590]=30'd858839683;
array2[18591]=30'd858839683;
array2[18592]=30'd865130113;
array2[18593]=30'd865130113;
array2[18594]=30'd858839683;
array2[18595]=30'd858839683;
array2[18596]=30'd858839683;
array2[18597]=30'd858839683;
array2[18598]=30'd858839683;
array2[18599]=30'd858839683;
array2[18600]=30'd858839683;
array2[18601]=30'd823228019;
array2[18602]=30'd319215128;
array2[18603]=30'd444954173;
array2[18604]=30'd858839683;
array2[18605]=30'd538207812;
array2[18606]=30'd193577377;
array2[18607]=30'd231362949;
array2[18608]=30'd234504581;
array2[18609]=30'd231362949;
array2[18610]=30'd230317442;
array2[18611]=30'd231362949;
array2[18612]=30'd229266819;
array2[18613]=30'd231362949;
array2[18614]=30'd234504581;
array2[18615]=30'd231362949;
array2[18616]=30'd231362949;
array2[18617]=30'd231362949;
array2[18618]=30'd229266819;
array2[18619]=30'd231362949;
array2[18620]=30'd231362949;
array2[18621]=30'd231362949;
array2[18622]=30'd234504581;
array2[18623]=30'd231362949;
array2[18624]=30'd823228019;
array2[18625]=30'd906004072;
array2[18626]=30'd906004072;
array2[18627]=30'd906004072;
array2[18628]=30'd736232864;
array2[18629]=30'd690121052;
array2[18630]=30'd690121052;
array2[18631]=30'd690121052;
array2[18632]=30'd690121052;
array2[18633]=30'd690121052;
array2[18634]=30'd690121052;
array2[18635]=30'd690121052;
array2[18636]=30'd690121052;
array2[18637]=30'd690121052;
array2[18638]=30'd690121052;
array2[18639]=30'd832648722;
array2[18640]=30'd906004072;
array2[18641]=30'd906004072;
array2[18642]=30'd906004072;
array2[18643]=30'd906004072;
array2[18644]=30'd906004072;
array2[18645]=30'd906004072;
array2[18646]=30'd906004072;
array2[18647]=30'd906004072;
array2[18648]=30'd906004072;
array2[18649]=30'd906004072;
array2[18650]=30'd906004072;
array2[18651]=30'd736232864;
array2[18652]=30'd690121052;
array2[18653]=30'd690121052;
array2[18654]=30'd690121052;
array2[18655]=30'd690121052;
array2[18656]=30'd690121052;
array2[18657]=30'd690121052;
array2[18658]=30'd690121052;
array2[18659]=30'd690121052;
array2[18660]=30'd690121052;
array2[18661]=30'd690121052;
array2[18662]=30'd281508345;
array2[18663]=30'd819020415;
array2[18664]=30'd851505800;
array2[18665]=30'd851505800;
array2[18666]=30'd851505800;
array2[18667]=30'd851505800;
array2[18668]=30'd858839683;
array2[18669]=30'd858839683;
array2[18670]=30'd858839683;
array2[18671]=30'd858839683;
array2[18672]=30'd858839683;
array2[18673]=30'd858839683;
array2[18674]=30'd858839683;
array2[18675]=30'd858839683;
array2[18676]=30'd858839683;
array2[18677]=30'd858839683;
array2[18678]=30'd858839683;
array2[18679]=30'd858839683;
array2[18680]=30'd865130113;
array2[18681]=30'd858839683;
array2[18682]=30'd865130113;
array2[18683]=30'd858839683;
array2[18684]=30'd865130113;
array2[18685]=30'd865130113;
array2[18686]=30'd865130113;
array2[18687]=30'd865130113;
array2[18688]=30'd858839683;
array2[18689]=30'd865130113;
array2[18690]=30'd858839683;
array2[18691]=30'd858839683;
array2[18692]=30'd858839683;
array2[18693]=30'd858839683;
array2[18694]=30'd865130113;
array2[18695]=30'd858839683;
array2[18696]=30'd858839683;
array2[18697]=30'd823228019;
array2[18698]=30'd347490866;
array2[18699]=30'd444954173;
array2[18700]=30'd819020415;
array2[18701]=30'd506770009;
array2[18702]=30'd193577377;
array2[18703]=30'd234504581;
array2[18704]=30'd234504581;
array2[18705]=30'd231362949;
array2[18706]=30'd231362949;
array2[18707]=30'd231362949;
array2[18708]=30'd230317442;
array2[18709]=30'd231364996;
array2[18710]=30'd234504581;
array2[18711]=30'd228216193;
array2[18712]=30'd231362949;
array2[18713]=30'd231362949;
array2[18714]=30'd230317442;
array2[18715]=30'd230317442;
array2[18716]=30'd231362949;
array2[18717]=30'd231362949;
array2[18718]=30'd231362949;
array2[18719]=30'd234504581;
array2[18720]=30'd639824186;
array2[18721]=30'd736232864;
array2[18722]=30'd690121052;
array2[18723]=30'd690121052;
array2[18724]=30'd637725975;
array2[18725]=30'd615715061;
array2[18726]=30'd615715061;
array2[18727]=30'd615715061;
array2[18728]=30'd611520752;
array2[18729]=30'd611520752;
array2[18730]=30'd611520752;
array2[18731]=30'd611520752;
array2[18732]=30'd611520752;
array2[18733]=30'd611520752;
array2[18734]=30'd611520752;
array2[18735]=30'd690121052;
array2[18736]=30'd690121052;
array2[18737]=30'd690121052;
array2[18738]=30'd690121052;
array2[18739]=30'd690121052;
array2[18740]=30'd736232864;
array2[18741]=30'd690121052;
array2[18742]=30'd690121052;
array2[18743]=30'd736232864;
array2[18744]=30'd736232864;
array2[18745]=30'd690121052;
array2[18746]=30'd736232864;
array2[18747]=30'd637725975;
array2[18748]=30'd611520752;
array2[18749]=30'd611520752;
array2[18750]=30'd611520752;
array2[18751]=30'd611520752;
array2[18752]=30'd611520752;
array2[18753]=30'd611520752;
array2[18754]=30'd611520752;
array2[18755]=30'd611520752;
array2[18756]=30'd606284005;
array2[18757]=30'd521469272;
array2[18758]=30'd352736774;
array2[18759]=30'd858839683;
array2[18760]=30'd865130113;
array2[18761]=30'd858839683;
array2[18762]=30'd858839683;
array2[18763]=30'd858839683;
array2[18764]=30'd865130113;
array2[18765]=30'd858839683;
array2[18766]=30'd858839683;
array2[18767]=30'd858839683;
array2[18768]=30'd858839683;
array2[18769]=30'd858839683;
array2[18770]=30'd858839683;
array2[18771]=30'd858839683;
array2[18772]=30'd858839683;
array2[18773]=30'd858839683;
array2[18774]=30'd858839683;
array2[18775]=30'd865130113;
array2[18776]=30'd865130113;
array2[18777]=30'd865130113;
array2[18778]=30'd865130113;
array2[18779]=30'd858839683;
array2[18780]=30'd858839683;
array2[18781]=30'd865130113;
array2[18782]=30'd858839683;
array2[18783]=30'd858839683;
array2[18784]=30'd858839683;
array2[18785]=30'd858839683;
array2[18786]=30'd865130113;
array2[18787]=30'd858839683;
array2[18788]=30'd858839683;
array2[18789]=30'd799112870;
array2[18790]=30'd732038833;
array2[18791]=30'd758240964;
array2[18792]=30'd851505800;
array2[18793]=30'd819020415;
array2[18794]=30'd434416250;
array2[18795]=30'd518272648;
array2[18796]=30'd828452495;
array2[18797]=30'd483727963;
array2[18798]=30'd179916222;
array2[18799]=30'd221916546;
array2[18800]=30'd227165569;
array2[18801]=30'd231362949;
array2[18802]=30'd231362949;
array2[18803]=30'd231362949;
array2[18804]=30'd229266819;
array2[18805]=30'd231362949;
array2[18806]=30'd234504581;
array2[18807]=30'd231362949;
array2[18808]=30'd231362949;
array2[18809]=30'd231362949;
array2[18810]=30'd231362949;
array2[18811]=30'd231362949;
array2[18812]=30'd231362949;
array2[18813]=30'd231362949;
array2[18814]=30'd234504581;
array2[18815]=30'd231359873;
array2[18816]=30'd582318295;
array2[18817]=30'd611520752;
array2[18818]=30'd615715061;
array2[18819]=30'd615715061;
array2[18820]=30'd615715061;
array2[18821]=30'd611520752;
array2[18822]=30'd606284005;
array2[18823]=30'd606284005;
array2[18824]=30'd606284005;
array2[18825]=30'd606284005;
array2[18826]=30'd606284005;
array2[18827]=30'd611520752;
array2[18828]=30'd611520752;
array2[18829]=30'd611520752;
array2[18830]=30'd611520752;
array2[18831]=30'd611520752;
array2[18832]=30'd611520752;
array2[18833]=30'd606284005;
array2[18834]=30'd606284005;
array2[18835]=30'd606284005;
array2[18836]=30'd606284005;
array2[18837]=30'd606284005;
array2[18838]=30'd611520752;
array2[18839]=30'd606284005;
array2[18840]=30'd606284005;
array2[18841]=30'd606284005;
array2[18842]=30'd606284005;
array2[18843]=30'd611520752;
array2[18844]=30'd611520752;
array2[18845]=30'd611520752;
array2[18846]=30'd611520752;
array2[18847]=30'd611520752;
array2[18848]=30'd611520752;
array2[18849]=30'd611520752;
array2[18850]=30'd611520752;
array2[18851]=30'd611520752;
array2[18852]=30'd611520752;
array2[18853]=30'd389419527;
array2[18854]=30'd483727963;
array2[18855]=30'd851505800;
array2[18856]=30'd865130113;
array2[18857]=30'd858839683;
array2[18858]=30'd858839683;
array2[18859]=30'd865130113;
array2[18860]=30'd865130113;
array2[18861]=30'd858839683;
array2[18862]=30'd858839683;
array2[18863]=30'd858839683;
array2[18864]=30'd858839683;
array2[18865]=30'd858839683;
array2[18866]=30'd858839683;
array2[18867]=30'd858839683;
array2[18868]=30'd858839683;
array2[18869]=30'd858839683;
array2[18870]=30'd865130113;
array2[18871]=30'd865130113;
array2[18872]=30'd865130113;
array2[18873]=30'd851505800;
array2[18874]=30'd858839683;
array2[18875]=30'd858839683;
array2[18876]=30'd858839683;
array2[18877]=30'd858839683;
array2[18878]=30'd858839683;
array2[18879]=30'd858839683;
array2[18880]=30'd858839683;
array2[18881]=30'd858839683;
array2[18882]=30'd865130113;
array2[18883]=30'd865130113;
array2[18884]=30'd770812573;
array2[18885]=30'd537140990;
array2[18886]=30'd409311115;
array2[18887]=30'd558174979;
array2[18888]=30'd758240964;
array2[18889]=30'd828452495;
array2[18890]=30'd677571193;
array2[18891]=30'd732038833;
array2[18892]=30'd828452495;
array2[18893]=30'd672348794;
array2[18894]=30'd299264555;
array2[18895]=30'd179916222;
array2[18896]=30'd232392085;
array2[18897]=30'd231359873;
array2[18898]=30'd234504581;
array2[18899]=30'd229266819;
array2[18900]=30'd231362949;
array2[18901]=30'd231362949;
array2[18902]=30'd231362949;
array2[18903]=30'd231362949;
array2[18904]=30'd231362949;
array2[18905]=30'd231362949;
array2[18906]=30'd228216193;
array2[18907]=30'd228216193;
array2[18908]=30'd229266819;
array2[18909]=30'd231362949;
array2[18910]=30'd230317442;
array2[18911]=30'd229266819;
array2[18912]=30'd582318295;
array2[18913]=30'd606284005;
array2[18914]=30'd611520752;
array2[18915]=30'd606284005;
array2[18916]=30'd585627858;
array2[18917]=30'd585627858;
array2[18918]=30'd585627858;
array2[18919]=30'd585627858;
array2[18920]=30'd585627858;
array2[18921]=30'd585627858;
array2[18922]=30'd585627858;
array2[18923]=30'd585627858;
array2[18924]=30'd585627858;
array2[18925]=30'd585627858;
array2[18926]=30'd585627858;
array2[18927]=30'd595854564;
array2[18928]=30'd615715061;
array2[18929]=30'd611520752;
array2[18930]=30'd611520752;
array2[18931]=30'd611520752;
array2[18932]=30'd611520752;
array2[18933]=30'd611520752;
array2[18934]=30'd611520752;
array2[18935]=30'd611520752;
array2[18936]=30'd611520752;
array2[18937]=30'd611520752;
array2[18938]=30'd611520752;
array2[18939]=30'd586531028;
array2[18940]=30'd585627858;
array2[18941]=30'd585627858;
array2[18942]=30'd585627858;
array2[18943]=30'd585627858;
array2[18944]=30'd585627858;
array2[18945]=30'd585627858;
array2[18946]=30'd585627858;
array2[18947]=30'd585627858;
array2[18948]=30'd585627858;
array2[18949]=30'd359161273;
array2[18950]=30'd678602388;
array2[18951]=30'd851505800;
array2[18952]=30'd865130113;
array2[18953]=30'd851505800;
array2[18954]=30'd851505800;
array2[18955]=30'd858839683;
array2[18956]=30'd858839683;
array2[18957]=30'd858839683;
array2[18958]=30'd858839683;
array2[18959]=30'd858839683;
array2[18960]=30'd858839683;
array2[18961]=30'd858839683;
array2[18962]=30'd858839683;
array2[18963]=30'd858839683;
array2[18964]=30'd858839683;
array2[18965]=30'd851505800;
array2[18966]=30'd858839683;
array2[18967]=30'd858839683;
array2[18968]=30'd858839683;
array2[18969]=30'd851505800;
array2[18970]=30'd858839683;
array2[18971]=30'd865130113;
array2[18972]=30'd865130113;
array2[18973]=30'd865130113;
array2[18974]=30'd858839683;
array2[18975]=30'd858839683;
array2[18976]=30'd865130113;
array2[18977]=30'd858839683;
array2[18978]=30'd858839683;
array2[18979]=30'd865130113;
array2[18980]=30'd539218630;
array2[18981]=30'd395649781;
array2[18982]=30'd390446940;
array2[18983]=30'd409311115;
array2[18984]=30'd558174979;
array2[18985]=30'd828452495;
array2[18986]=30'd858839683;
array2[18987]=30'd851505800;
array2[18988]=30'd858839683;
array2[18989]=30'd828452495;
array2[18990]=30'd678602388;
array2[18991]=30'd265736724;
array2[18992]=30'd220861839;
array2[18993]=30'd231362949;
array2[18994]=30'd231362949;
array2[18995]=30'd229266819;
array2[18996]=30'd231362949;
array2[18997]=30'd234504581;
array2[18998]=30'd229266819;
array2[18999]=30'd231362949;
array2[19000]=30'd234504581;
array2[19001]=30'd227165569;
array2[19002]=30'd231362949;
array2[19003]=30'd231362949;
array2[19004]=30'd231362949;
array2[19005]=30'd229266819;
array2[19006]=30'd231362949;
array2[19007]=30'd229266819;
array2[19008]=30'd561572038;
array2[19009]=30'd561572038;
array2[19010]=30'd561572038;
array2[19011]=30'd561572038;
array2[19012]=30'd514590904;
array2[19013]=30'd524037312;
array2[19014]=30'd518815920;
array2[19015]=30'd518815920;
array2[19016]=30'd518815920;
array2[19017]=30'd518815920;
array2[19018]=30'd518815920;
array2[19019]=30'd518815920;
array2[19020]=30'd518815920;
array2[19021]=30'd518815920;
array2[19022]=30'd524037312;
array2[19023]=30'd543866052;
array2[19024]=30'd561572038;
array2[19025]=30'd561572038;
array2[19026]=30'd561572038;
array2[19027]=30'd561572038;
array2[19028]=30'd561572038;
array2[19029]=30'd561572038;
array2[19030]=30'd561572038;
array2[19031]=30'd561572038;
array2[19032]=30'd561572038;
array2[19033]=30'd561572038;
array2[19034]=30'd561572038;
array2[19035]=30'd514590904;
array2[19036]=30'd518815920;
array2[19037]=30'd518815920;
array2[19038]=30'd518815920;
array2[19039]=30'd518815920;
array2[19040]=30'd518815920;
array2[19041]=30'd518815920;
array2[19042]=30'd518815920;
array2[19043]=30'd518815920;
array2[19044]=30'd518815920;
array2[19045]=30'd338288022;
array2[19046]=30'd711090860;
array2[19047]=30'd851505800;
array2[19048]=30'd851505800;
array2[19049]=30'd858839683;
array2[19050]=30'd865130113;
array2[19051]=30'd865130113;
array2[19052]=30'd858839683;
array2[19053]=30'd858839683;
array2[19054]=30'd851505800;
array2[19055]=30'd828452495;
array2[19056]=30'd851505800;
array2[19057]=30'd828452495;
array2[19058]=30'd770812573;
array2[19059]=30'd770812573;
array2[19060]=30'd770812573;
array2[19061]=30'd758240964;
array2[19062]=30'd799112870;
array2[19063]=30'd858839683;
array2[19064]=30'd858839683;
array2[19065]=30'd865130113;
array2[19066]=30'd858839683;
array2[19067]=30'd865130113;
array2[19068]=30'd865130113;
array2[19069]=30'd858839683;
array2[19070]=30'd858839683;
array2[19071]=30'd858839683;
array2[19072]=30'd858839683;
array2[19073]=30'd858839683;
array2[19074]=30'd858839683;
array2[19075]=30'd851505800;
array2[19076]=30'd395649781;
array2[19077]=30'd395649781;
array2[19078]=30'd451191548;
array2[19079]=30'd390446940;
array2[19080]=30'd409311115;
array2[19081]=30'd770812573;
array2[19082]=30'd851505800;
array2[19083]=30'd851505800;
array2[19084]=30'd851505800;
array2[19085]=30'd828452495;
array2[19086]=30'd764529268;
array2[19087]=30'd319215128;
array2[19088]=30'd232392085;
array2[19089]=30'd231362949;
array2[19090]=30'd231362949;
array2[19091]=30'd231362949;
array2[19092]=30'd231362949;
array2[19093]=30'd231362949;
array2[19094]=30'd231362949;
array2[19095]=30'd231362949;
array2[19096]=30'd231362949;
array2[19097]=30'd231362949;
array2[19098]=30'd231362949;
array2[19099]=30'd231359873;
array2[19100]=30'd230317442;
array2[19101]=30'd229266819;
array2[19102]=30'd231362949;
array2[19103]=30'd231362949;
array2[19104]=30'd530274492;
array2[19105]=30'd521966763;
array2[19106]=30'd521966763;
array2[19107]=30'd521966763;
array2[19108]=30'd521966763;
array2[19109]=30'd521966763;
array2[19110]=30'd521966763;
array2[19111]=30'd521966763;
array2[19112]=30'd521966763;
array2[19113]=30'd521966763;
array2[19114]=30'd521966763;
array2[19115]=30'd521966763;
array2[19116]=30'd521966763;
array2[19117]=30'd521966763;
array2[19118]=30'd521966763;
array2[19119]=30'd521966763;
array2[19120]=30'd521966763;
array2[19121]=30'd521966763;
array2[19122]=30'd518815920;
array2[19123]=30'd521966763;
array2[19124]=30'd521966763;
array2[19125]=30'd521966763;
array2[19126]=30'd521966763;
array2[19127]=30'd518815920;
array2[19128]=30'd518815920;
array2[19129]=30'd521966763;
array2[19130]=30'd521966763;
array2[19131]=30'd521966763;
array2[19132]=30'd521966763;
array2[19133]=30'd521966763;
array2[19134]=30'd521966763;
array2[19135]=30'd521966763;
array2[19136]=30'd521966763;
array2[19137]=30'd521966763;
array2[19138]=30'd521966763;
array2[19139]=30'd521966763;
array2[19140]=30'd521966763;
array2[19141]=30'd301610387;
array2[19142]=30'd711090860;
array2[19143]=30'd851505800;
array2[19144]=30'd858839683;
array2[19145]=30'd858839683;
array2[19146]=30'd858839683;
array2[19147]=30'd858839683;
array2[19148]=30'd828452495;
array2[19149]=30'd799112870;
array2[19150]=30'd672348794;
array2[19151]=30'd678602388;
array2[19152]=30'd770812573;
array2[19153]=30'd770812573;
array2[19154]=30'd732038833;
array2[19155]=30'd732038833;
array2[19156]=30'd732038833;
array2[19157]=30'd732038833;
array2[19158]=30'd732038833;
array2[19159]=30'd770812573;
array2[19160]=30'd770812573;
array2[19161]=30'd851505800;
array2[19162]=30'd858839683;
array2[19163]=30'd858839683;
array2[19164]=30'd851505800;
array2[19165]=30'd858839683;
array2[19166]=30'd865130113;
array2[19167]=30'd865130113;
array2[19168]=30'd865130113;
array2[19169]=30'd858839683;
array2[19170]=30'd858839683;
array2[19171]=30'd858839683;
array2[19172]=30'd732038833;
array2[19173]=30'd451191548;
array2[19174]=30'd451191548;
array2[19175]=30'd451191548;
array2[19176]=30'd713202349;
array2[19177]=30'd828452495;
array2[19178]=30'd851505800;
array2[19179]=30'd858839683;
array2[19180]=30'd858839683;
array2[19181]=30'd727851632;
array2[19182]=30'd401997362;
array2[19183]=30'd228181405;
array2[19184]=30'd227165569;
array2[19185]=30'd230317442;
array2[19186]=30'd231362949;
array2[19187]=30'd229266819;
array2[19188]=30'd231362949;
array2[19189]=30'd231362949;
array2[19190]=30'd231362949;
array2[19191]=30'd230317442;
array2[19192]=30'd231362949;
array2[19193]=30'd231362949;
array2[19194]=30'd228216193;
array2[19195]=30'd231362949;
array2[19196]=30'd231362949;
array2[19197]=30'd231362949;
array2[19198]=30'd231362949;
array2[19199]=30'd227165569;
array2[19200]=30'd530274492;
array2[19201]=30'd521966763;
array2[19202]=30'd521966763;
array2[19203]=30'd521966763;
array2[19204]=30'd515671261;
array2[19205]=30'd510427417;
array2[19206]=30'd510427417;
array2[19207]=30'd510427417;
array2[19208]=30'd510427417;
array2[19209]=30'd510427417;
array2[19210]=30'd510427417;
array2[19211]=30'd510427417;
array2[19212]=30'd510427417;
array2[19213]=30'd510427417;
array2[19214]=30'd510427417;
array2[19215]=30'd839470532;
array2[19216]=30'd777593273;
array2[19217]=30'd521966763;
array2[19218]=30'd521966763;
array2[19219]=30'd521966763;
array2[19220]=30'd521966763;
array2[19221]=30'd521966763;
array2[19222]=30'd521966763;
array2[19223]=30'd521966763;
array2[19224]=30'd521966763;
array2[19225]=30'd521966763;
array2[19226]=30'd521966763;
array2[19227]=30'd515671261;
array2[19228]=30'd510427417;
array2[19229]=30'd510427417;
array2[19230]=30'd510427417;
array2[19231]=30'd510427417;
array2[19232]=30'd510427417;
array2[19233]=30'd510427417;
array2[19234]=30'd510427417;
array2[19235]=30'd510427417;
array2[19236]=30'd496710898;
array2[19237]=30'd381167075;
array2[19238]=30'd764529268;
array2[19239]=30'd764529268;
array2[19240]=30'd799112870;
array2[19241]=30'd828452495;
array2[19242]=30'd828452495;
array2[19243]=30'd799112870;
array2[19244]=30'd732038833;
array2[19245]=30'd678602388;
array2[19246]=30'd450208341;
array2[19247]=30'd560184961;
array2[19248]=30'd606320275;
array2[19249]=30'd631447172;
array2[19250]=30'd631447172;
array2[19251]=30'd606320275;
array2[19252]=30'd631447172;
array2[19253]=30'd678602388;
array2[19254]=30'd732038833;
array2[19255]=30'd732038833;
array2[19256]=30'd732038833;
array2[19257]=30'd770812573;
array2[19258]=30'd851505800;
array2[19259]=30'd858839683;
array2[19260]=30'd851505800;
array2[19261]=30'd851505800;
array2[19262]=30'd858839683;
array2[19263]=30'd858839683;
array2[19264]=30'd851505800;
array2[19265]=30'd828452495;
array2[19266]=30'd858839683;
array2[19267]=30'd858839683;
array2[19268]=30'd858839683;
array2[19269]=30'd758240964;
array2[19270]=30'd582196031;
array2[19271]=30'd672324351;
array2[19272]=30'd828452495;
array2[19273]=30'd851505800;
array2[19274]=30'd858839683;
array2[19275]=30'd858839683;
array2[19276]=30'd828452495;
array2[19277]=30'd762499681;
array2[19278]=30'd383147560;
array2[19279]=30'd232392085;
array2[19280]=30'd227165569;
array2[19281]=30'd231364996;
array2[19282]=30'd231364996;
array2[19283]=30'd231364996;
array2[19284]=30'd230317442;
array2[19285]=30'd229266819;
array2[19286]=30'd231359873;
array2[19287]=30'd230317442;
array2[19288]=30'd231362949;
array2[19289]=30'd230317442;
array2[19290]=30'd231362949;
array2[19291]=30'd231362949;
array2[19292]=30'd230317442;
array2[19293]=30'd229266819;
array2[19294]=30'd231359873;
array2[19295]=30'd228216193;
array2[19296]=30'd462205301;
array2[19297]=30'd482131304;
array2[19298]=30'd482131304;
array2[19299]=30'd475838865;
array2[19300]=30'd477946350;
array2[19301]=30'd482138634;
array2[19302]=30'd475850257;
array2[19303]=30'd482138634;
array2[19304]=30'd482138634;
array2[19305]=30'd482138634;
array2[19306]=30'd475850257;
array2[19307]=30'd482138634;
array2[19308]=30'd475850257;
array2[19309]=30'd482138634;
array2[19310]=30'd473746934;
array2[19311]=30'd608913932;
array2[19312]=30'd608913932;
array2[19313]=30'd482131304;
array2[19314]=30'd482131304;
array2[19315]=30'd482131304;
array2[19316]=30'd482131304;
array2[19317]=30'd482131304;
array2[19318]=30'd482131304;
array2[19319]=30'd482131304;
array2[19320]=30'd482131304;
array2[19321]=30'd482131304;
array2[19322]=30'd482131304;
array2[19323]=30'd473746934;
array2[19324]=30'd482138634;
array2[19325]=30'd482138634;
array2[19326]=30'd482138634;
array2[19327]=30'd482138634;
array2[19328]=30'd482138634;
array2[19329]=30'd482138634;
array2[19330]=30'd475850257;
array2[19331]=30'd482138634;
array2[19332]=30'd307963313;
array2[19333]=30'd631447172;
array2[19334]=30'd805398138;
array2[19335]=30'd407216718;
array2[19336]=30'd606320275;
array2[19337]=30'd631447172;
array2[19338]=30'd606320275;
array2[19339]=30'd560184961;
array2[19340]=30'd560184961;
array2[19341]=30'd434416250;
array2[19342]=30'd302686639;
array2[19343]=30'd307963313;
array2[19344]=30'd207191473;
array2[19345]=30'd179916222;
array2[19346]=30'd179916222;
array2[19347]=30'd179916222;
array2[19348]=30'd179916222;
array2[19349]=30'd347490866;
array2[19350]=30'd566515308;
array2[19351]=30'd560184961;
array2[19352]=30'd678602388;
array2[19353]=30'd711090860;
array2[19354]=30'd711090860;
array2[19355]=30'd828452495;
array2[19356]=30'd851505800;
array2[19357]=30'd858839683;
array2[19358]=30'd858839683;
array2[19359]=30'd858839683;
array2[19360]=30'd805398138;
array2[19361]=30'd711090860;
array2[19362]=30'd799112870;
array2[19363]=30'd828452495;
array2[19364]=30'd851505800;
array2[19365]=30'd858839683;
array2[19366]=30'd858839683;
array2[19367]=30'd851505800;
array2[19368]=30'd851505800;
array2[19369]=30'd851505800;
array2[19370]=30'd828452495;
array2[19371]=30'd828452495;
array2[19372]=30'd678602388;
array2[19373]=30'd401997362;
array2[19374]=30'd212454818;
array2[19375]=30'd227165569;
array2[19376]=30'd231359873;
array2[19377]=30'd231362949;
array2[19378]=30'd231362949;
array2[19379]=30'd231364996;
array2[19380]=30'd231362949;
array2[19381]=30'd229270912;
array2[19382]=30'd231362949;
array2[19383]=30'd231362949;
array2[19384]=30'd227165569;
array2[19385]=30'd230317442;
array2[19386]=30'd231362949;
array2[19387]=30'd231362949;
array2[19388]=30'd230317442;
array2[19389]=30'd231362949;
array2[19390]=30'd229266819;
array2[19391]=30'd231362949;
array2[19392]=30'd457992679;
array2[19393]=30'd475850257;
array2[19394]=30'd482138634;
array2[19395]=30'd475850257;
array2[19396]=30'd480046615;
array2[19397]=30'd475850257;
array2[19398]=30'd480046615;
array2[19399]=30'd475850257;
array2[19400]=30'd480046615;
array2[19401]=30'd475850257;
array2[19402]=30'd475850257;
array2[19403]=30'd480046615;
array2[19404]=30'd482138634;
array2[19405]=30'd480046615;
array2[19406]=30'd480046615;
array2[19407]=30'd480046615;
array2[19408]=30'd480046615;
array2[19409]=30'd475850257;
array2[19410]=30'd482138634;
array2[19411]=30'd480046615;
array2[19412]=30'd475850257;
array2[19413]=30'd480046615;
array2[19414]=30'd480046615;
array2[19415]=30'd480046615;
array2[19416]=30'd475850257;
array2[19417]=30'd480046615;
array2[19418]=30'd482138634;
array2[19419]=30'd480046615;
array2[19420]=30'd475850257;
array2[19421]=30'd480046615;
array2[19422]=30'd480046615;
array2[19423]=30'd475850257;
array2[19424]=30'd480046615;
array2[19425]=30'd475850257;
array2[19426]=30'd475850257;
array2[19427]=30'd480046615;
array2[19428]=30'd302686639;
array2[19429]=30'd631447172;
array2[19430]=30'd483727963;
array2[19431]=30'd178773498;
array2[19432]=30'd304706973;
array2[19433]=30'd387723742;
array2[19434]=30'd340509129;
array2[19435]=30'd340509129;
array2[19436]=30'd340509129;
array2[19437]=30'd387723742;
array2[19438]=30'd475850257;
array2[19439]=30'd490515973;
array2[19440]=30'd307963313;
array2[19441]=30'd228216193;
array2[19442]=30'd230317442;
array2[19443]=30'd229270912;
array2[19444]=30'd229270912;
array2[19445]=30'd232392085;
array2[19446]=30'd193577377;
array2[19447]=30'd193577377;
array2[19448]=30'd347490866;
array2[19449]=30'd357913199;
array2[19450]=30'd606320275;
array2[19451]=30'd732038833;
array2[19452]=30'd828452495;
array2[19453]=30'd858839683;
array2[19454]=30'd858839683;
array2[19455]=30'd858839683;
array2[19456]=30'd764529268;
array2[19457]=30'd631447172;
array2[19458]=30'd770812573;
array2[19459]=30'd732038833;
array2[19460]=30'd770812573;
array2[19461]=30'd799112870;
array2[19462]=30'd799112870;
array2[19463]=30'd799112870;
array2[19464]=30'd770812573;
array2[19465]=30'd770812573;
array2[19466]=30'd604201637;
array2[19467]=30'd407216718;
array2[19468]=30'd319215128;
array2[19469]=30'd213516691;
array2[19470]=30'd234504581;
array2[19471]=30'd228216193;
array2[19472]=30'd231359873;
array2[19473]=30'd231359873;
array2[19474]=30'd231362949;
array2[19475]=30'd231362949;
array2[19476]=30'd231362949;
array2[19477]=30'd234504581;
array2[19478]=30'd227165569;
array2[19479]=30'd231362949;
array2[19480]=30'd231362949;
array2[19481]=30'd231362949;
array2[19482]=30'd228216193;
array2[19483]=30'd229266819;
array2[19484]=30'd231362949;
array2[19485]=30'd227165569;
array2[19486]=30'd230317442;
array2[19487]=30'd229266819;
array2[19488]=30'd439121402;
array2[19489]=30'd475850257;
array2[19490]=30'd475850257;
array2[19491]=30'd482138634;
array2[19492]=30'd457992679;
array2[19493]=30'd439121402;
array2[19494]=30'd439121402;
array2[19495]=30'd439121402;
array2[19496]=30'd387723742;
array2[19497]=30'd439121402;
array2[19498]=30'd387723742;
array2[19499]=30'd816426489;
array2[19500]=30'd608913932;
array2[19501]=30'd439121402;
array2[19502]=30'd439121402;
array2[19503]=30'd473746934;
array2[19504]=30'd482138634;
array2[19505]=30'd480046615;
array2[19506]=30'd475850257;
array2[19507]=30'd608913932;
array2[19508]=30'd608913932;
array2[19509]=30'd490515973;
array2[19510]=30'd475850257;
array2[19511]=30'd482138634;
array2[19512]=30'd480046615;
array2[19513]=30'd475850257;
array2[19514]=30'd475850257;
array2[19515]=30'd457992679;
array2[19516]=30'd439121402;
array2[19517]=30'd439121402;
array2[19518]=30'd439121402;
array2[19519]=30'd439121402;
array2[19520]=30'd439121402;
array2[19521]=30'd439121402;
array2[19522]=30'd608913932;
array2[19523]=30'd608913932;
array2[19524]=30'd232434043;
array2[19525]=30'd347490866;
array2[19526]=30'd362496490;
array2[19527]=30'd150539724;
array2[19528]=30'd302686639;
array2[19529]=30'd480046615;
array2[19530]=30'd608913932;
array2[19531]=30'd816426489;
array2[19532]=30'd490515973;
array2[19533]=30'd480046615;
array2[19534]=30'd475850257;
array2[19535]=30'd473746934;
array2[19536]=30'd302686639;
array2[19537]=30'd231362949;
array2[19538]=30'd229266819;
array2[19539]=30'd227165569;
array2[19540]=30'd228216193;
array2[19541]=30'd231364996;
array2[19542]=30'd231362949;
array2[19543]=30'd228216193;
array2[19544]=30'd212454818;
array2[19545]=30'd207191473;
array2[19546]=30'd450208341;
array2[19547]=30'd711090860;
array2[19548]=30'd799112870;
array2[19549]=30'd858839683;
array2[19550]=30'd851505800;
array2[19551]=30'd865130113;
array2[19552]=30'd764529268;
array2[19553]=30'd560184961;
array2[19554]=30'd711090860;
array2[19555]=30'd732038833;
array2[19556]=30'd732038833;
array2[19557]=30'd732038833;
array2[19558]=30'd732038833;
array2[19559]=30'd732038833;
array2[19560]=30'd678602388;
array2[19561]=30'd450208341;
array2[19562]=30'd319215128;
array2[19563]=30'd212454818;
array2[19564]=30'd213516691;
array2[19565]=30'd234504581;
array2[19566]=30'd228216193;
array2[19567]=30'd231362949;
array2[19568]=30'd234504581;
array2[19569]=30'd229266819;
array2[19570]=30'd229270912;
array2[19571]=30'd231362949;
array2[19572]=30'd230317442;
array2[19573]=30'd230317442;
array2[19574]=30'd229266819;
array2[19575]=30'd228216193;
array2[19576]=30'd231359873;
array2[19577]=30'd230317442;
array2[19578]=30'd230317442;
array2[19579]=30'd229270912;
array2[19580]=30'd230317442;
array2[19581]=30'd231362949;
array2[19582]=30'd230317442;
array2[19583]=30'd231362949;
array2[19584]=30'd340509129;
array2[19585]=30'd387723742;
array2[19586]=30'd387723742;
array2[19587]=30'd340509129;
array2[19588]=30'd265985428;
array2[19589]=30'd229270912;
array2[19590]=30'd229270912;
array2[19591]=30'd229266819;
array2[19592]=30'd229266819;
array2[19593]=30'd228212100;
array2[19594]=30'd238691720;
array2[19595]=30'd719920570;
array2[19596]=30'd616102353;
array2[19597]=30'd227159434;
array2[19598]=30'd234515845;
array2[19599]=30'd340509129;
array2[19600]=30'd387723742;
array2[19601]=30'd387723742;
array2[19602]=30'd387723742;
array2[19603]=30'd719920570;
array2[19604]=30'd719920570;
array2[19605]=30'd340509129;
array2[19606]=30'd387723742;
array2[19607]=30'd387723742;
array2[19608]=30'd387723742;
array2[19609]=30'd387723742;
array2[19610]=30'd387723742;
array2[19611]=30'd302686639;
array2[19612]=30'd229270912;
array2[19613]=30'd229270912;
array2[19614]=30'd231364996;
array2[19615]=30'd225072515;
array2[19616]=30'd229266819;
array2[19617]=30'd231362949;
array2[19618]=30'd664345022;
array2[19619]=30'd670611929;
array2[19620]=30'd248105365;
array2[19621]=30'd213516691;
array2[19622]=30'd307963313;
array2[19623]=30'd307963313;
array2[19624]=30'd362496490;
array2[19625]=30'd387723742;
array2[19626]=30'd655981997;
array2[19627]=30'd747191732;
array2[19628]=30'd362496490;
array2[19629]=30'd387723742;
array2[19630]=30'd387723742;
array2[19631]=30'd340509129;
array2[19632]=30'd265985428;
array2[19633]=30'd231364996;
array2[19634]=30'd231364996;
array2[19635]=30'd230317442;
array2[19636]=30'd230317442;
array2[19637]=30'd228216193;
array2[19638]=30'd229266819;
array2[19639]=30'd231362949;
array2[19640]=30'd229266819;
array2[19641]=30'd228216193;
array2[19642]=30'd260631016;
array2[19643]=30'd518272648;
array2[19644]=30'd732038833;
array2[19645]=30'd828452495;
array2[19646]=30'd858839683;
array2[19647]=30'd851505800;
array2[19648]=30'd819020415;
array2[19649]=30'd560184961;
array2[19650]=30'd518272648;
array2[19651]=30'd518272648;
array2[19652]=30'd518272648;
array2[19653]=30'd483727963;
array2[19654]=30'd319215128;
array2[19655]=30'd319215128;
array2[19656]=30'd319215128;
array2[19657]=30'd212454818;
array2[19658]=30'd221916546;
array2[19659]=30'd230317442;
array2[19660]=30'd231362949;
array2[19661]=30'd230317442;
array2[19662]=30'd231362949;
array2[19663]=30'd228216193;
array2[19664]=30'd231362949;
array2[19665]=30'd231364996;
array2[19666]=30'd230317442;
array2[19667]=30'd229270912;
array2[19668]=30'd230317442;
array2[19669]=30'd231362949;
array2[19670]=30'd231362949;
array2[19671]=30'd231362949;
array2[19672]=30'd234504581;
array2[19673]=30'd228216193;
array2[19674]=30'd231362949;
array2[19675]=30'd231362949;
array2[19676]=30'd231362949;
array2[19677]=30'd230317442;
array2[19678]=30'd231362949;
array2[19679]=30'd231362949;
array2[19680]=30'd212454818;
array2[19681]=30'd234504581;
array2[19682]=30'd236604812;
array2[19683]=30'd229270912;
array2[19684]=30'd231364996;
array2[19685]=30'd231364996;
array2[19686]=30'd231362949;
array2[19687]=30'd234504581;
array2[19688]=30'd231362949;
array2[19689]=30'd231359873;
array2[19690]=30'd231362949;
array2[19691]=30'd231364996;
array2[19692]=30'd225072515;
array2[19693]=30'd231362949;
array2[19694]=30'd231362949;
array2[19695]=30'd230317442;
array2[19696]=30'd227165569;
array2[19697]=30'd228216193;
array2[19698]=30'd227165569;
array2[19699]=30'd227165569;
array2[19700]=30'd227159434;
array2[19701]=30'd231362949;
array2[19702]=30'd227165569;
array2[19703]=30'd231362949;
array2[19704]=30'd227165569;
array2[19705]=30'd227165569;
array2[19706]=30'd228216193;
array2[19707]=30'd229266819;
array2[19708]=30'd230317442;
array2[19709]=30'd229266819;
array2[19710]=30'd230317442;
array2[19711]=30'd229266819;
array2[19712]=30'd231362949;
array2[19713]=30'd231364996;
array2[19714]=30'd231362949;
array2[19715]=30'd231359873;
array2[19716]=30'd227165569;
array2[19717]=30'd231362949;
array2[19718]=30'd231362949;
array2[19719]=30'd227165569;
array2[19720]=30'd227165569;
array2[19721]=30'd228216193;
array2[19722]=30'd225072515;
array2[19723]=30'd227165569;
array2[19724]=30'd231362949;
array2[19725]=30'd227165569;
array2[19726]=30'd227165569;
array2[19727]=30'd231362949;
array2[19728]=30'd227165569;
array2[19729]=30'd231364996;
array2[19730]=30'd231364996;
array2[19731]=30'd231362949;
array2[19732]=30'd229266819;
array2[19733]=30'd231362949;
array2[19734]=30'd229266819;
array2[19735]=30'd231362949;
array2[19736]=30'd230317442;
array2[19737]=30'd231362949;
array2[19738]=30'd186252693;
array2[19739]=30'd407216718;
array2[19740]=30'd678602388;
array2[19741]=30'd770812573;
array2[19742]=30'd851505800;
array2[19743]=30'd858839683;
array2[19744]=30'd858839683;
array2[19745]=30'd646130287;
array2[19746]=30'd481587821;
array2[19747]=30'd539218630;
array2[19748]=30'd485780117;
array2[19749]=30'd190356956;
array2[19750]=30'd221916546;
array2[19751]=30'd231362949;
array2[19752]=30'd225072515;
array2[19753]=30'd229270912;
array2[19754]=30'd231362949;
array2[19755]=30'd230317442;
array2[19756]=30'd231362949;
array2[19757]=30'd231364996;
array2[19758]=30'd231362949;
array2[19759]=30'd229266819;
array2[19760]=30'd228216193;
array2[19761]=30'd229266819;
array2[19762]=30'd231364996;
array2[19763]=30'd230317442;
array2[19764]=30'd230317442;
array2[19765]=30'd229266819;
array2[19766]=30'd231362949;
array2[19767]=30'd231362949;
array2[19768]=30'd234504581;
array2[19769]=30'd231362949;
array2[19770]=30'd228216193;
array2[19771]=30'd231362949;
array2[19772]=30'd231362949;
array2[19773]=30'd229266819;
array2[19774]=30'd230317442;
array2[19775]=30'd229266819;
array2[19776]=30'd228181405;
array2[19777]=30'd227165569;
array2[19778]=30'd228216193;
array2[19779]=30'd232417668;
array2[19780]=30'd231364996;
array2[19781]=30'd231364996;
array2[19782]=30'd231362949;
array2[19783]=30'd231362949;
array2[19784]=30'd228216193;
array2[19785]=30'd234504581;
array2[19786]=30'd231362949;
array2[19787]=30'd231362949;
array2[19788]=30'd231362949;
array2[19789]=30'd231362949;
array2[19790]=30'd234504581;
array2[19791]=30'd532258209;
array2[19792]=30'd532258209;
array2[19793]=30'd228212100;
array2[19794]=30'd231362949;
array2[19795]=30'd229266819;
array2[19796]=30'd230317442;
array2[19797]=30'd229266819;
array2[19798]=30'd231362949;
array2[19799]=30'd231359873;
array2[19800]=30'd231362949;
array2[19801]=30'd231362949;
array2[19802]=30'd229266819;
array2[19803]=30'd231362949;
array2[19804]=30'd231362949;
array2[19805]=30'd227165569;
array2[19806]=30'd231362949;
array2[19807]=30'd231362949;
array2[19808]=30'd234504581;
array2[19809]=30'd228216193;
array2[19810]=30'd231362949;
array2[19811]=30'd234504581;
array2[19812]=30'd231362949;
array2[19813]=30'd225072515;
array2[19814]=30'd472496545;
array2[19815]=30'd616102353;
array2[19816]=30'd238691720;
array2[19817]=30'd231362949;
array2[19818]=30'd230317442;
array2[19819]=30'd230317442;
array2[19820]=30'd231362949;
array2[19821]=30'd228216193;
array2[19822]=30'd229266819;
array2[19823]=30'd231362949;
array2[19824]=30'd231362949;
array2[19825]=30'd231362949;
array2[19826]=30'd231364996;
array2[19827]=30'd234504581;
array2[19828]=30'd231362949;
array2[19829]=30'd231362949;
array2[19830]=30'd231362949;
array2[19831]=30'd231362949;
array2[19832]=30'd229266819;
array2[19833]=30'd229266819;
array2[19834]=30'd228216193;
array2[19835]=30'd212454818;
array2[19836]=30'd407216718;
array2[19837]=30'd678602388;
array2[19838]=30'd770812573;
array2[19839]=30'd851505800;
array2[19840]=30'd858839683;
array2[19841]=30'd708987491;
array2[19842]=30'd485780117;
array2[19843]=30'd606320275;
array2[19844]=30'd539218630;
array2[19845]=30'd299264555;
array2[19846]=30'd220861839;
array2[19847]=30'd231362949;
array2[19848]=30'd229270912;
array2[19849]=30'd229266819;
array2[19850]=30'd231364996;
array2[19851]=30'd231362949;
array2[19852]=30'd231362949;
array2[19853]=30'd230317442;
array2[19854]=30'd231362949;
array2[19855]=30'd230317442;
array2[19856]=30'd231362949;
array2[19857]=30'd231362949;
array2[19858]=30'd231362949;
array2[19859]=30'd231362949;
array2[19860]=30'd231362949;
array2[19861]=30'd231362949;
array2[19862]=30'd231362949;
array2[19863]=30'd231362949;
array2[19864]=30'd231362949;
array2[19865]=30'd230317442;
array2[19866]=30'd229266819;
array2[19867]=30'd231362949;
array2[19868]=30'd229266819;
array2[19869]=30'd231362949;
array2[19870]=30'd231364996;
array2[19871]=30'd229266819;
array2[19872]=30'd212454818;
array2[19873]=30'd234504581;
array2[19874]=30'd228212100;
array2[19875]=30'd231359873;
array2[19876]=30'd231362949;
array2[19877]=30'd231362949;
array2[19878]=30'd227165569;
array2[19879]=30'd234504581;
array2[19880]=30'd231359873;
array2[19881]=30'd231362949;
array2[19882]=30'd231362949;
array2[19883]=30'd231362949;
array2[19884]=30'd231362949;
array2[19885]=30'd231359873;
array2[19886]=30'd256519562;
array2[19887]=30'd719920570;
array2[19888]=30'd664345022;
array2[19889]=30'd210373000;
array2[19890]=30'd234504581;
array2[19891]=30'd227165569;
array2[19892]=30'd230317442;
array2[19893]=30'd231364996;
array2[19894]=30'd231362949;
array2[19895]=30'd229266819;
array2[19896]=30'd231362949;
array2[19897]=30'd230317442;
array2[19898]=30'd231362949;
array2[19899]=30'd231364996;
array2[19900]=30'd231362949;
array2[19901]=30'd234504581;
array2[19902]=30'd231362949;
array2[19903]=30'd231362949;
array2[19904]=30'd231362949;
array2[19905]=30'd231362949;
array2[19906]=30'd231362949;
array2[19907]=30'd231362949;
array2[19908]=30'd229266819;
array2[19909]=30'd228212100;
array2[19910]=30'd616102353;
array2[19911]=30'd777593273;
array2[19912]=30'd238691720;
array2[19913]=30'd231362949;
array2[19914]=30'd231362949;
array2[19915]=30'd229270912;
array2[19916]=30'd231362949;
array2[19917]=30'd229266819;
array2[19918]=30'd229266819;
array2[19919]=30'd229266819;
array2[19920]=30'd231362949;
array2[19921]=30'd231364996;
array2[19922]=30'd229270912;
array2[19923]=30'd231362949;
array2[19924]=30'd231362949;
array2[19925]=30'd227165569;
array2[19926]=30'd230317442;
array2[19927]=30'd234504581;
array2[19928]=30'd231362949;
array2[19929]=30'd231364996;
array2[19930]=30'd229266819;
array2[19931]=30'd229266819;
array2[19932]=30'd195647926;
array2[19933]=30'd606320275;
array2[19934]=30'd732038833;
array2[19935]=30'd828452495;
array2[19936]=30'd858839683;
array2[19937]=30'd828452495;
array2[19938]=30'd560184961;
array2[19939]=30'd539218630;
array2[19940]=30'd601041592;
array2[19941]=30'd485780117;
array2[19942]=30'd179916222;
array2[19943]=30'd230317442;
array2[19944]=30'd231362949;
array2[19945]=30'd231362949;
array2[19946]=30'd229266819;
array2[19947]=30'd231362949;
array2[19948]=30'd231362949;
array2[19949]=30'd231362949;
array2[19950]=30'd231362949;
array2[19951]=30'd231362949;
array2[19952]=30'd234504581;
array2[19953]=30'd231362949;
array2[19954]=30'd231362949;
array2[19955]=30'd231362949;
array2[19956]=30'd231362949;
array2[19957]=30'd231362949;
array2[19958]=30'd234504581;
array2[19959]=30'd231362949;
array2[19960]=30'd231362949;
array2[19961]=30'd231362949;
array2[19962]=30'd229266819;
array2[19963]=30'd229266819;
array2[19964]=30'd230317442;
array2[19965]=30'd229266819;
array2[19966]=30'd234504581;
array2[19967]=30'd228216193;
array2[19968]=30'd212454818;
array2[19969]=30'd234504581;
array2[19970]=30'd228212100;
array2[19971]=30'd229266819;
array2[19972]=30'd234504581;
array2[19973]=30'd231362949;
array2[19974]=30'd227165569;
array2[19975]=30'd231362949;
array2[19976]=30'd228216193;
array2[19977]=30'd234504581;
array2[19978]=30'd231362949;
array2[19979]=30'd231362949;
array2[19980]=30'd231362949;
array2[19981]=30'd231362949;
array2[19982]=30'd227165569;
array2[19983]=30'd231362949;
array2[19984]=30'd236604812;
array2[19985]=30'd231362949;
array2[19986]=30'd229270912;
array2[19987]=30'd231362949;
array2[19988]=30'd230317442;
array2[19989]=30'd234504581;
array2[19990]=30'd231362949;
array2[19991]=30'd229266819;
array2[19992]=30'd229266819;
array2[19993]=30'd229266819;
array2[19994]=30'd231359873;
array2[19995]=30'd231362949;
array2[19996]=30'd231362949;
array2[19997]=30'd231359873;
array2[19998]=30'd234504581;
array2[19999]=30'd228216193;
array2[20000]=30'd231362949;
array2[20001]=30'd231362949;
array2[20002]=30'd231362949;
array2[20003]=30'd231362949;
array2[20004]=30'd229266819;
array2[20005]=30'd234504581;
array2[20006]=30'd236604812;
array2[20007]=30'd231364996;
array2[20008]=30'd231364996;
array2[20009]=30'd228212100;
array2[20010]=30'd230317442;
array2[20011]=30'd232417668;
array2[20012]=30'd231362949;
array2[20013]=30'd229266819;
array2[20014]=30'd231362949;
array2[20015]=30'd229266819;
array2[20016]=30'd231362949;
array2[20017]=30'd231362949;
array2[20018]=30'd234504581;
array2[20019]=30'd231362949;
array2[20020]=30'd231362949;
array2[20021]=30'd228216193;
array2[20022]=30'd230317442;
array2[20023]=30'd234504581;
array2[20024]=30'd229266819;
array2[20025]=30'd234504581;
array2[20026]=30'd231364996;
array2[20027]=30'd231362949;
array2[20028]=30'd212454818;
array2[20029]=30'd407216718;
array2[20030]=30'd601041592;
array2[20031]=30'd770812573;
array2[20032]=30'd851505800;
array2[20033]=30'd858839683;
array2[20034]=30'd565444213;
array2[20035]=30'd539218630;
array2[20036]=30'd601041592;
array2[20037]=30'd539218630;
array2[20038]=30'd295074390;
array2[20039]=30'd213516691;
array2[20040]=30'd231359873;
array2[20041]=30'd231364996;
array2[20042]=30'd229266819;
array2[20043]=30'd229266819;
array2[20044]=30'd228216193;
array2[20045]=30'd228216193;
array2[20046]=30'd231362949;
array2[20047]=30'd231362949;
array2[20048]=30'd231364996;
array2[20049]=30'd231362949;
array2[20050]=30'd231362949;
array2[20051]=30'd231362949;
array2[20052]=30'd228216193;
array2[20053]=30'd231362949;
array2[20054]=30'd234504581;
array2[20055]=30'd231362949;
array2[20056]=30'd231362949;
array2[20057]=30'd229266819;
array2[20058]=30'd229266819;
array2[20059]=30'd229266819;
array2[20060]=30'd231362949;
array2[20061]=30'd231364996;
array2[20062]=30'd234504581;
array2[20063]=30'd231362949;
array2[20064]=30'd228181405;
array2[20065]=30'd234504581;
array2[20066]=30'd227159434;
array2[20067]=30'd231359873;
array2[20068]=30'd231362949;
array2[20069]=30'd231362949;
array2[20070]=30'd230307208;
array2[20071]=30'd234504581;
array2[20072]=30'd234504581;
array2[20073]=30'd228216193;
array2[20074]=30'd231359873;
array2[20075]=30'd231362949;
array2[20076]=30'd231362949;
array2[20077]=30'd231362949;
array2[20078]=30'd231362949;
array2[20079]=30'd234504581;
array2[20080]=30'd231362949;
array2[20081]=30'd231359873;
array2[20082]=30'd231362949;
array2[20083]=30'd229266819;
array2[20084]=30'd229266819;
array2[20085]=30'd230317442;
array2[20086]=30'd231362949;
array2[20087]=30'd234504581;
array2[20088]=30'd229266819;
array2[20089]=30'd229266819;
array2[20090]=30'd228216193;
array2[20091]=30'd231362949;
array2[20092]=30'd231362949;
array2[20093]=30'd231364996;
array2[20094]=30'd231362949;
array2[20095]=30'd229266819;
array2[20096]=30'd234504581;
array2[20097]=30'd231362949;
array2[20098]=30'd231362949;
array2[20099]=30'd231362949;
array2[20100]=30'd231362949;
array2[20101]=30'd231362949;
array2[20102]=30'd231359873;
array2[20103]=30'd231364996;
array2[20104]=30'd229266819;
array2[20105]=30'd231362949;
array2[20106]=30'd229266819;
array2[20107]=30'd231362949;
array2[20108]=30'd234504581;
array2[20109]=30'd234504581;
array2[20110]=30'd234504581;
array2[20111]=30'd231362949;
array2[20112]=30'd231362949;
array2[20113]=30'd230317442;
array2[20114]=30'd230317442;
array2[20115]=30'd229266819;
array2[20116]=30'd231362949;
array2[20117]=30'd231359873;
array2[20118]=30'd231364996;
array2[20119]=30'd231359873;
array2[20120]=30'd231362949;
array2[20121]=30'd231364996;
array2[20122]=30'd231364996;
array2[20123]=30'd229266819;
array2[20124]=30'd230317442;
array2[20125]=30'd228181405;
array2[20126]=30'd338018898;
array2[20127]=30'd711090860;
array2[20128]=30'd770812573;
array2[20129]=30'd828452495;
array2[20130]=30'd606320275;
array2[20131]=30'd518272648;
array2[20132]=30'd539218630;
array2[20133]=30'd601041592;
array2[20134]=30'd434416250;
array2[20135]=30'd195647926;
array2[20136]=30'd228216193;
array2[20137]=30'd229270912;
array2[20138]=30'd229266819;
array2[20139]=30'd229266819;
array2[20140]=30'd231359873;
array2[20141]=30'd228216193;
array2[20142]=30'd231362949;
array2[20143]=30'd231362949;
array2[20144]=30'd231362949;
array2[20145]=30'd234504581;
array2[20146]=30'd230317442;
array2[20147]=30'd230317442;
array2[20148]=30'd229266819;
array2[20149]=30'd231362949;
array2[20150]=30'd231364996;
array2[20151]=30'd231362949;
array2[20152]=30'd229266819;
array2[20153]=30'd231359873;
array2[20154]=30'd231362949;
array2[20155]=30'd229266819;
array2[20156]=30'd230317442;
array2[20157]=30'd231364996;
array2[20158]=30'd231364996;
array2[20159]=30'd230317442;
array2[20160]=30'd212454818;
array2[20161]=30'd234504581;
array2[20162]=30'd228212100;
array2[20163]=30'd229266819;
array2[20164]=30'd234504581;
array2[20165]=30'd231362949;
array2[20166]=30'd227165569;
array2[20167]=30'd231362949;
array2[20168]=30'd234504581;
array2[20169]=30'd234504581;
array2[20170]=30'd231362949;
array2[20171]=30'd231362949;
array2[20172]=30'd231362949;
array2[20173]=30'd231362949;
array2[20174]=30'd229266819;
array2[20175]=30'd231362949;
array2[20176]=30'd231362949;
array2[20177]=30'd231362949;
array2[20178]=30'd231359873;
array2[20179]=30'd231362949;
array2[20180]=30'd230317442;
array2[20181]=30'd230317442;
array2[20182]=30'd230317442;
array2[20183]=30'd231362949;
array2[20184]=30'd231362949;
array2[20185]=30'd229266819;
array2[20186]=30'd231362949;
array2[20187]=30'd227165569;
array2[20188]=30'd231364996;
array2[20189]=30'd231362949;
array2[20190]=30'd231362949;
array2[20191]=30'd229266819;
array2[20192]=30'd230317442;
array2[20193]=30'd234504581;
array2[20194]=30'd231362949;
array2[20195]=30'd234504581;
array2[20196]=30'd231362949;
array2[20197]=30'd231364996;
array2[20198]=30'd228212100;
array2[20199]=30'd231364996;
array2[20200]=30'd231362949;
array2[20201]=30'd231362949;
array2[20202]=30'd231362949;
array2[20203]=30'd229266819;
array2[20204]=30'd229266819;
array2[20205]=30'd231362949;
array2[20206]=30'd231362949;
array2[20207]=30'd231362949;
array2[20208]=30'd231362949;
array2[20209]=30'd231362949;
array2[20210]=30'd229266819;
array2[20211]=30'd229266819;
array2[20212]=30'd230317442;
array2[20213]=30'd230317442;
array2[20214]=30'd231362949;
array2[20215]=30'd234504581;
array2[20216]=30'd231362949;
array2[20217]=30'd229266819;
array2[20218]=30'd228216193;
array2[20219]=30'd228216193;
array2[20220]=30'd231364996;
array2[20221]=30'd227159434;
array2[20222]=30'd190356956;
array2[20223]=30'd606320275;
array2[20224]=30'd732038833;
array2[20225]=30'd770812573;
array2[20226]=30'd713179821;
array2[20227]=30'd347490866;
array2[20228]=30'd299264555;
array2[20229]=30'd518272648;
array2[20230]=30'd518272648;
array2[20231]=30'd347490866;
array2[20232]=30'd220861839;
array2[20233]=30'd231364996;
array2[20234]=30'd229266819;
array2[20235]=30'd229266819;
array2[20236]=30'd230317442;
array2[20237]=30'd229266819;
array2[20238]=30'd229266819;
array2[20239]=30'd228216193;
array2[20240]=30'd231362949;
array2[20241]=30'd231362949;
array2[20242]=30'd231364996;
array2[20243]=30'd234504581;
array2[20244]=30'd231362949;
array2[20245]=30'd231364996;
array2[20246]=30'd229266819;
array2[20247]=30'd231362949;
array2[20248]=30'd228216193;
array2[20249]=30'd229266819;
array2[20250]=30'd234504581;
array2[20251]=30'd231362949;
array2[20252]=30'd231362949;
array2[20253]=30'd229266819;
array2[20254]=30'd231362949;
array2[20255]=30'd230317442;
array2[20256]=30'd212454818;
array2[20257]=30'd234504581;
array2[20258]=30'd228212100;
array2[20259]=30'd231362949;
array2[20260]=30'd234504581;
array2[20261]=30'd231362949;
array2[20262]=30'd228216193;
array2[20263]=30'd230317442;
array2[20264]=30'd231362949;
array2[20265]=30'd234504581;
array2[20266]=30'd229266819;
array2[20267]=30'd231362949;
array2[20268]=30'd231362949;
array2[20269]=30'd231362949;
array2[20270]=30'd228216193;
array2[20271]=30'd231362949;
array2[20272]=30'd231362949;
array2[20273]=30'd229266819;
array2[20274]=30'd231359873;
array2[20275]=30'd231362949;
array2[20276]=30'd231362949;
array2[20277]=30'd229266819;
array2[20278]=30'd231364996;
array2[20279]=30'd228216193;
array2[20280]=30'd231362949;
array2[20281]=30'd231364996;
array2[20282]=30'd231362949;
array2[20283]=30'd228216193;
array2[20284]=30'd228216193;
array2[20285]=30'd231362949;
array2[20286]=30'd234504581;
array2[20287]=30'd228216193;
array2[20288]=30'd231362949;
array2[20289]=30'd231362949;
array2[20290]=30'd231362949;
array2[20291]=30'd231362949;
array2[20292]=30'd231362949;
array2[20293]=30'd231362949;
array2[20294]=30'd231362949;
array2[20295]=30'd227165569;
array2[20296]=30'd231362949;
array2[20297]=30'd231362949;
array2[20298]=30'd229266819;
array2[20299]=30'd231362949;
array2[20300]=30'd229266819;
array2[20301]=30'd230317442;
array2[20302]=30'd231362949;
array2[20303]=30'd231362949;
array2[20304]=30'd231359873;
array2[20305]=30'd231362949;
array2[20306]=30'd228216193;
array2[20307]=30'd231362949;
array2[20308]=30'd231362949;
array2[20309]=30'd231362949;
array2[20310]=30'd231359873;
array2[20311]=30'd231362949;
array2[20312]=30'd234504581;
array2[20313]=30'd231362949;
array2[20314]=30'd231362949;
array2[20315]=30'd231362949;
array2[20316]=30'd230317442;
array2[20317]=30'd231362949;
array2[20318]=30'd220861839;
array2[20319]=30'd383147560;
array2[20320]=30'd606320275;
array2[20321]=30'd678602388;
array2[20322]=30'd631447172;
array2[20323]=30'd299264555;
array2[20324]=30'd254365107;
array2[20325]=30'd401997362;
array2[20326]=30'd319215128;
array2[20327]=30'd319215128;
array2[20328]=30'd213516691;
array2[20329]=30'd227165569;
array2[20330]=30'd229266819;
array2[20331]=30'd231362949;
array2[20332]=30'd231362949;
array2[20333]=30'd231362949;
array2[20334]=30'd229266819;
array2[20335]=30'd231362949;
array2[20336]=30'd229266819;
array2[20337]=30'd231362949;
array2[20338]=30'd231362949;
array2[20339]=30'd231362949;
array2[20340]=30'd231362949;
array2[20341]=30'd231362949;
array2[20342]=30'd229266819;
array2[20343]=30'd229266819;
array2[20344]=30'd231362949;
array2[20345]=30'd231362949;
array2[20346]=30'd234504581;
array2[20347]=30'd231362949;
array2[20348]=30'd231362949;
array2[20349]=30'd228216193;
array2[20350]=30'd230317442;
array2[20351]=30'd231362949;
array2[20352]=30'd212454818;
array2[20353]=30'd234504581;
array2[20354]=30'd228212100;
array2[20355]=30'd229266819;
array2[20356]=30'd234504581;
array2[20357]=30'd231362949;
array2[20358]=30'd227165569;
array2[20359]=30'd231362949;
array2[20360]=30'd234504581;
array2[20361]=30'd234504581;
array2[20362]=30'd230317442;
array2[20363]=30'd229266819;
array2[20364]=30'd228216193;
array2[20365]=30'd231362949;
array2[20366]=30'd231362949;
array2[20367]=30'd230317442;
array2[20368]=30'd230317442;
array2[20369]=30'd230317442;
array2[20370]=30'd231362949;
array2[20371]=30'd231362949;
array2[20372]=30'd231362949;
array2[20373]=30'd231362949;
array2[20374]=30'd231362949;
array2[20375]=30'd231364996;
array2[20376]=30'd231362949;
array2[20377]=30'd231362949;
array2[20378]=30'd229266819;
array2[20379]=30'd229266819;
array2[20380]=30'd234504581;
array2[20381]=30'd231362949;
array2[20382]=30'd231362949;
array2[20383]=30'd231362949;
array2[20384]=30'd230317442;
array2[20385]=30'd228216193;
array2[20386]=30'd228216193;
array2[20387]=30'd231362949;
array2[20388]=30'd229266819;
array2[20389]=30'd231362949;
array2[20390]=30'd230317442;
array2[20391]=30'd228216193;
array2[20392]=30'd227165569;
array2[20393]=30'd230317442;
array2[20394]=30'd231362949;
array2[20395]=30'd231364996;
array2[20396]=30'd229266819;
array2[20397]=30'd231362949;
array2[20398]=30'd229266819;
array2[20399]=30'd231362949;
array2[20400]=30'd231362949;
array2[20401]=30'd230317442;
array2[20402]=30'd229270912;
array2[20403]=30'd229266819;
array2[20404]=30'd229266819;
array2[20405]=30'd229266819;
array2[20406]=30'd231362949;
array2[20407]=30'd234504581;
array2[20408]=30'd231362949;
array2[20409]=30'd234504581;
array2[20410]=30'd231362949;
array2[20411]=30'd229266819;
array2[20412]=30'd230317442;
array2[20413]=30'd231362949;
array2[20414]=30'd231362949;
array2[20415]=30'd213516691;
array2[20416]=30'd281508345;
array2[20417]=30'd281508345;
array2[20418]=30'd319215128;
array2[20419]=30'd190356956;
array2[20420]=30'd232392085;
array2[20421]=30'd238691720;
array2[20422]=30'd234499470;
array2[20423]=30'd238691720;
array2[20424]=30'd231362949;
array2[20425]=30'd231362949;
array2[20426]=30'd230317442;
array2[20427]=30'd231362949;
array2[20428]=30'd231362949;
array2[20429]=30'd228216193;
array2[20430]=30'd230317442;
array2[20431]=30'd230317442;
array2[20432]=30'd231362949;
array2[20433]=30'd231362949;
array2[20434]=30'd231364996;
array2[20435]=30'd230317442;
array2[20436]=30'd229266819;
array2[20437]=30'd234504581;
array2[20438]=30'd231362949;
array2[20439]=30'd231362949;
array2[20440]=30'd231362949;
array2[20441]=30'd231362949;
array2[20442]=30'd231362949;
array2[20443]=30'd231362949;
array2[20444]=30'd231362949;
array2[20445]=30'd229266819;
array2[20446]=30'd231362949;
array2[20447]=30'd231364996;
array2[20448]=30'd212454818;
array2[20449]=30'd231359873;
array2[20450]=30'd227165569;
array2[20451]=30'd231362949;
array2[20452]=30'd234504581;
array2[20453]=30'd231362949;
array2[20454]=30'd231362949;
array2[20455]=30'd230317442;
array2[20456]=30'd231362949;
array2[20457]=30'd234504581;
array2[20458]=30'd230317442;
array2[20459]=30'd229266819;
array2[20460]=30'd231362949;
array2[20461]=30'd231362949;
array2[20462]=30'd228216193;
array2[20463]=30'd230317442;
array2[20464]=30'd230317442;
array2[20465]=30'd231362949;
array2[20466]=30'd229266819;
array2[20467]=30'd231362949;
array2[20468]=30'd228216193;
array2[20469]=30'd231364996;
array2[20470]=30'd230317442;
array2[20471]=30'd231364996;
array2[20472]=30'd230317442;
array2[20473]=30'd228216193;
array2[20474]=30'd231364996;
array2[20475]=30'd231362949;
array2[20476]=30'd234504581;
array2[20477]=30'd228216193;
array2[20478]=30'd231364996;
array2[20479]=30'd231362949;
array2[20480]=30'd229266819;
array2[20481]=30'd231362949;
array2[20482]=30'd230317442;
array2[20483]=30'd231362949;
array2[20484]=30'd231362949;
array2[20485]=30'd231359873;
array2[20486]=30'd230317442;
array2[20487]=30'd231364996;
array2[20488]=30'd227159434;
array2[20489]=30'd231364996;
array2[20490]=30'd231362949;
array2[20491]=30'd231362949;
array2[20492]=30'd229266819;
array2[20493]=30'd229266819;
array2[20494]=30'd231362949;
array2[20495]=30'd229266819;
array2[20496]=30'd231362949;
array2[20497]=30'd231362949;
array2[20498]=30'd231362949;
array2[20499]=30'd231364996;
array2[20500]=30'd229266819;
array2[20501]=30'd230317442;
array2[20502]=30'd231362949;
array2[20503]=30'd229266819;
array2[20504]=30'd231362949;
array2[20505]=30'd234504581;
array2[20506]=30'd231362949;
array2[20507]=30'd231362949;
array2[20508]=30'd229266819;
array2[20509]=30'd231362949;
array2[20510]=30'd231362949;
array2[20511]=30'd231362949;
array2[20512]=30'd227165569;
array2[20513]=30'd227165569;
array2[20514]=30'd227165569;
array2[20515]=30'd230307208;
array2[20516]=30'd231362949;
array2[20517]=30'd231362949;
array2[20518]=30'd231362949;
array2[20519]=30'd230317442;
array2[20520]=30'd231362949;
array2[20521]=30'd231362949;
array2[20522]=30'd231362949;
array2[20523]=30'd229266819;
array2[20524]=30'd231362949;
array2[20525]=30'd231362949;
array2[20526]=30'd231364996;
array2[20527]=30'd230317442;
array2[20528]=30'd231359873;
array2[20529]=30'd231362949;
array2[20530]=30'd228216193;
array2[20531]=30'd231362949;
array2[20532]=30'd231362949;
array2[20533]=30'd231362949;
array2[20534]=30'd228216193;
array2[20535]=30'd231362949;
array2[20536]=30'd231362949;
array2[20537]=30'd231362949;
array2[20538]=30'd234504581;
array2[20539]=30'd231362949;
array2[20540]=30'd231362949;
array2[20541]=30'd230317442;
array2[20542]=30'd231362949;
array2[20543]=30'd228212100;
array2[20544]=30'd212454818;
array2[20545]=30'd234504581;
array2[20546]=30'd228212100;
array2[20547]=30'd229266819;
array2[20548]=30'd234504581;
array2[20549]=30'd231362949;
array2[20550]=30'd227165569;
array2[20551]=30'd231362949;
array2[20552]=30'd234504581;
array2[20553]=30'd234504581;
array2[20554]=30'd229266819;
array2[20555]=30'd229266819;
array2[20556]=30'd231362949;
array2[20557]=30'd231362949;
array2[20558]=30'd228216193;
array2[20559]=30'd229266819;
array2[20560]=30'd229266819;
array2[20561]=30'd234504581;
array2[20562]=30'd227165569;
array2[20563]=30'd231362949;
array2[20564]=30'd231362949;
array2[20565]=30'd231362949;
array2[20566]=30'd231362949;
array2[20567]=30'd231362949;
array2[20568]=30'd231359873;
array2[20569]=30'd234504581;
array2[20570]=30'd228216193;
array2[20571]=30'd231362949;
array2[20572]=30'd231362949;
array2[20573]=30'd231362949;
array2[20574]=30'd231362949;
array2[20575]=30'd231362949;
array2[20576]=30'd234504581;
array2[20577]=30'd231362949;
array2[20578]=30'd231362949;
array2[20579]=30'd234504581;
array2[20580]=30'd231362949;
array2[20581]=30'd234504581;
array2[20582]=30'd231364996;
array2[20583]=30'd231362949;
array2[20584]=30'd229266819;
array2[20585]=30'd231362949;
array2[20586]=30'd231362949;
array2[20587]=30'd234504581;
array2[20588]=30'd231362949;
array2[20589]=30'd231362949;
array2[20590]=30'd231362949;
array2[20591]=30'd231362949;
array2[20592]=30'd231362949;
array2[20593]=30'd231362949;
array2[20594]=30'd234504581;
array2[20595]=30'd229266819;
array2[20596]=30'd234504581;
array2[20597]=30'd231362949;
array2[20598]=30'd231362949;
array2[20599]=30'd231362949;
array2[20600]=30'd231362949;
array2[20601]=30'd234504581;
array2[20602]=30'd231362949;
array2[20603]=30'd231359873;
array2[20604]=30'd231364996;
array2[20605]=30'd231364996;
array2[20606]=30'd230317442;
array2[20607]=30'd229266819;
array2[20608]=30'd231362949;
array2[20609]=30'd231362949;
array2[20610]=30'd231359873;
array2[20611]=30'd227165569;
array2[20612]=30'd228216193;
array2[20613]=30'd231362949;
array2[20614]=30'd231364996;
array2[20615]=30'd231362949;
array2[20616]=30'd231362949;
array2[20617]=30'd231362949;
array2[20618]=30'd231359873;
array2[20619]=30'd231362949;
array2[20620]=30'd231362949;
array2[20621]=30'd231362949;
array2[20622]=30'd230317442;
array2[20623]=30'd231362949;
array2[20624]=30'd231362949;
array2[20625]=30'd234504581;
array2[20626]=30'd231362949;
array2[20627]=30'd231364996;
array2[20628]=30'd231362949;
array2[20629]=30'd229266819;
array2[20630]=30'd231362949;
array2[20631]=30'd234504581;
array2[20632]=30'd231359873;
array2[20633]=30'd231362949;
array2[20634]=30'd231362949;
array2[20635]=30'd231362949;
array2[20636]=30'd229266819;
array2[20637]=30'd230317442;
array2[20638]=30'd229266819;
array2[20639]=30'd234504581;
array2[20640]=30'd212454818;
array2[20641]=30'd231359873;
array2[20642]=30'd228216193;
array2[20643]=30'd234504581;
array2[20644]=30'd234504581;
array2[20645]=30'd231362949;
array2[20646]=30'd231362949;
array2[20647]=30'd229266819;
array2[20648]=30'd231362949;
array2[20649]=30'd234504581;
array2[20650]=30'd231362949;
array2[20651]=30'd231362949;
array2[20652]=30'd231359873;
array2[20653]=30'd231364996;
array2[20654]=30'd229266819;
array2[20655]=30'd230317442;
array2[20656]=30'd230317442;
array2[20657]=30'd231362949;
array2[20658]=30'd231362949;
array2[20659]=30'd229266819;
array2[20660]=30'd231362949;
array2[20661]=30'd228216193;
array2[20662]=30'd231362949;
array2[20663]=30'd231364996;
array2[20664]=30'd231362949;
array2[20665]=30'd230317442;
array2[20666]=30'd229266819;
array2[20667]=30'd234504581;
array2[20668]=30'd230317442;
array2[20669]=30'd234504581;
array2[20670]=30'd234504581;
array2[20671]=30'd231362949;
array2[20672]=30'd231362949;
array2[20673]=30'd231362949;
array2[20674]=30'd231362949;
array2[20675]=30'd231362949;
array2[20676]=30'd230317442;
array2[20677]=30'd231362949;
array2[20678]=30'd229266819;
array2[20679]=30'd231362949;
array2[20680]=30'd230317442;
array2[20681]=30'd234504581;
array2[20682]=30'd227165569;
array2[20683]=30'd230317442;
array2[20684]=30'd230317442;
array2[20685]=30'd229266819;
array2[20686]=30'd231362949;
array2[20687]=30'd229266819;
array2[20688]=30'd231362949;
array2[20689]=30'd228216193;
array2[20690]=30'd231362949;
array2[20691]=30'd229266819;
array2[20692]=30'd234504581;
array2[20693]=30'd231362949;
array2[20694]=30'd231362949;
array2[20695]=30'd231362949;
array2[20696]=30'd231362949;
array2[20697]=30'd231362949;
array2[20698]=30'd231362949;
array2[20699]=30'd231362949;
array2[20700]=30'd227165569;
array2[20701]=30'd228216193;
array2[20702]=30'd230317442;
array2[20703]=30'd229266819;
array2[20704]=30'd229266819;
array2[20705]=30'd229266819;
array2[20706]=30'd229266819;
array2[20707]=30'd231362949;
array2[20708]=30'd229266819;
array2[20709]=30'd231362949;
array2[20710]=30'd228216193;
array2[20711]=30'd231362949;
array2[20712]=30'd231364996;
array2[20713]=30'd231362949;
array2[20714]=30'd229266819;
array2[20715]=30'd229266819;
array2[20716]=30'd231362949;
array2[20717]=30'd231362949;
array2[20718]=30'd231362949;
array2[20719]=30'd231362949;
array2[20720]=30'd231362949;
array2[20721]=30'd231362949;
array2[20722]=30'd231364996;
array2[20723]=30'd231362949;
array2[20724]=30'd234504581;
array2[20725]=30'd230317442;
array2[20726]=30'd231364996;
array2[20727]=30'd229266819;
array2[20728]=30'd228216193;
array2[20729]=30'd229266819;
array2[20730]=30'd229266819;
array2[20731]=30'd230317442;
array2[20732]=30'd230317442;
array2[20733]=30'd230317442;
array2[20734]=30'd231362949;
array2[20735]=30'd272255371;



array[0]=30'd856066696;
array[1]=30'd856066696;
array[2]=30'd856066696;
array[3]=30'd856066696;
array[4]=30'd856066696;
array[5]=30'd856066696;
array[6]=30'd856066696;
array[7]=30'd856066696;
array[8]=30'd856066696;
array[9]=30'd856066696;
array[10]=30'd856066696;
array[11]=30'd856066696;
array[12]=30'd856066696;
array[13]=30'd856066696;
array[14]=30'd856066696;
array[15]=30'd856066696;
array[16]=30'd856066696;
array[17]=30'd856066696;
array[18]=30'd856066696;
array[19]=30'd856066696;
array[20]=30'd856066696;
array[21]=30'd856066696;
array[22]=30'd856066696;
array[23]=30'd856066696;
array[24]=30'd856066696;
array[25]=30'd856066696;
array[26]=30'd856066696;
array[27]=30'd856066696;
array[28]=30'd879168118;
array[29]=30'd884420162;
array[30]=30'd860309028;
array[31]=30'd843548160;
array[32]=30'd903304711;
array[33]=30'd810005031;
array[34]=30'd860309028;
array[35]=30'd841408084;
array[36]=30'd856066696;
array[37]=30'd856066696;
array[38]=30'd856066696;
array[39]=30'd856066696;
array[40]=30'd856066696;
array[41]=30'd856066696;
array[42]=30'd856066696;
array[43]=30'd729186945;
array[44]=30'd467006094;
array[45]=30'd496374434;
array[46]=30'd559255224;
array[47]=30'd608527024;
array[48]=30'd608527024;
array[49]=30'd547692230;
array[50]=30'd633661142;
array[51]=30'd633661142;
array[52]=30'd581260986;
array[53]=30'd581260986;
array[54]=30'd650433234;
array[55]=30'd633661142;
array[56]=30'd608527024;
array[57]=30'd653676161;
array[58]=30'd522581659;
array[59]=30'd646262454;
array[60]=30'd650433234;
array[61]=30'd633661142;
array[62]=30'd633661142;
array[63]=30'd650433234;
array[64]=30'd650433234;
array[65]=30'd650433234;
array[66]=30'd633661142;
array[67]=30'd633661142;
array[68]=30'd650433234;
array[69]=30'd581260986;
array[70]=30'd362130088;
array[71]=30'd581260986;
array[72]=30'd646262454;
array[73]=30'd633661142;
array[74]=30'd633661142;
array[75]=30'd633661142;
array[76]=30'd633661142;
array[77]=30'd650433234;
array[78]=30'd633661142;
array[79]=30'd613805729;
array[80]=30'd814111379;
array[81]=30'd824623759;
array[82]=30'd824623759;
array[83]=30'd824623759;
array[84]=30'd824623759;
array[85]=30'd856066696;
array[86]=30'd856066696;
array[87]=30'd824623759;
array[88]=30'd856066696;
array[89]=30'd856066696;
array[90]=30'd856066696;
array[91]=30'd856066696;
array[92]=30'd856066696;
array[93]=30'd856066696;
array[94]=30'd856066696;
array[95]=30'd824623759;
array[96]=30'd856066696;
array[97]=30'd856066696;
array[98]=30'd856066696;
array[99]=30'd856066696;
array[100]=30'd856066696;
array[101]=30'd856066696;
array[102]=30'd856066696;
array[103]=30'd856066696;
array[104]=30'd856066696;
array[105]=30'd856066696;
array[106]=30'd856066696;
array[107]=30'd856066696;
array[108]=30'd856066696;
array[109]=30'd856066696;
array[110]=30'd856066696;
array[111]=30'd856066696;
array[112]=30'd856066696;
array[113]=30'd856066696;
array[114]=30'd856066696;
array[115]=30'd856066696;
array[116]=30'd856066696;
array[117]=30'd856066696;
array[118]=30'd856066696;
array[119]=30'd856066696;
array[120]=30'd856066696;
array[121]=30'd856066696;
array[122]=30'd856066696;
array[123]=30'd856066696;
array[124]=30'd879168118;
array[125]=30'd879168118;
array[126]=30'd884420162;
array[127]=30'd860309028;
array[128]=30'd860309028;
array[129]=30'd841408084;
array[130]=30'd841408084;
array[131]=30'd856066696;
array[132]=30'd856066696;
array[133]=30'd856066696;
array[134]=30'd856066696;
array[135]=30'd856066696;
array[136]=30'd856066696;
array[137]=30'd856066696;
array[138]=30'd824623759;
array[139]=30'd582343294;
array[140]=30'd452327079;
array[141]=30'd613805729;
array[142]=30'd444952244;
array[143]=30'd646262454;
array[144]=30'd516257448;
array[145]=30'd608527024;
array[146]=30'd646262454;
array[147]=30'd646262454;
array[148]=30'd516257448;
array[149]=30'd633661142;
array[150]=30'd650433234;
array[151]=30'd646262454;
array[152]=30'd551919254;
array[153]=30'd815194717;
array[154]=30'd527847013;
array[155]=30'd608527024;
array[156]=30'd633661142;
array[157]=30'd633661142;
array[158]=30'd633661142;
array[159]=30'd633661142;
array[160]=30'd650433234;
array[161]=30'd650433234;
array[162]=30'd633661142;
array[163]=30'd633661142;
array[164]=30'd633661142;
array[165]=30'd646262454;
array[166]=30'd427157133;
array[167]=30'd496374434;
array[168]=30'd646262454;
array[169]=30'd633661142;
array[170]=30'd633661142;
array[171]=30'd633661142;
array[172]=30'd646262454;
array[173]=30'd633661142;
array[174]=30'd633661142;
array[175]=30'd581260986;
array[176]=30'd725995173;
array[177]=30'd824623759;
array[178]=30'd856066696;
array[179]=30'd856066696;
array[180]=30'd856066696;
array[181]=30'd814111379;
array[182]=30'd856066696;
array[183]=30'd856066696;
array[184]=30'd856066696;
array[185]=30'd856066696;
array[186]=30'd856066696;
array[187]=30'd856066696;
array[188]=30'd856066696;
array[189]=30'd856066696;
array[190]=30'd856066696;
array[191]=30'd879168118;
array[192]=30'd856066696;
array[193]=30'd856066696;
array[194]=30'd856066696;
array[195]=30'd856066696;
array[196]=30'd856066696;
array[197]=30'd856066696;
array[198]=30'd856066696;
array[199]=30'd856066696;
array[200]=30'd729186945;
array[201]=30'd709306968;
array[202]=30'd824623759;
array[203]=30'd856066696;
array[204]=30'd856066696;
array[205]=30'd856066696;
array[206]=30'd856066696;
array[207]=30'd856066696;
array[208]=30'd856066696;
array[209]=30'd856066696;
array[210]=30'd856066696;
array[211]=30'd856066696;
array[212]=30'd856066696;
array[213]=30'd856066696;
array[214]=30'd856066696;
array[215]=30'd856066696;
array[216]=30'd856066696;
array[217]=30'd856066696;
array[218]=30'd856066696;
array[219]=30'd856066696;
array[220]=30'd856066696;
array[221]=30'd856066696;
array[222]=30'd879168118;
array[223]=30'd841408084;
array[224]=30'd841408084;
array[225]=30'd841408084;
array[226]=30'd856066696;
array[227]=30'd856066696;
array[228]=30'd856066696;
array[229]=30'd856066696;
array[230]=30'd856066696;
array[231]=30'd856066696;
array[232]=30'd856066696;
array[233]=30'd856066696;
array[234]=30'd781608573;
array[235]=30'd496374434;
array[236]=30'd467006094;
array[237]=30'd634745492;
array[238]=30'd485848753;
array[239]=30'd646262454;
array[240]=30'd485848753;
array[241]=30'd646262454;
array[242]=30'd646262454;
array[243]=30'd646262454;
array[244]=30'd516257448;
array[245]=30'd646262454;
array[246]=30'd650433234;
array[247]=30'd559255224;
array[248]=30'd739680847;
array[249]=30'd815194717;
array[250]=30'd527847013;
array[251]=30'd608527024;
array[252]=30'd633661142;
array[253]=30'd633661142;
array[254]=30'd633661142;
array[255]=30'd633661142;
array[256]=30'd633661142;
array[257]=30'd650433234;
array[258]=30'd633661142;
array[259]=30'd633661142;
array[260]=30'd633661142;
array[261]=30'd633661142;
array[262]=30'd485848753;
array[263]=30'd362130088;
array[264]=30'd646262454;
array[265]=30'd633661142;
array[266]=30'd633661142;
array[267]=30'd633661142;
array[268]=30'd547692230;
array[269]=30'd608527024;
array[270]=30'd633661142;
array[271]=30'd646262454;
array[272]=30'd551919254;
array[273]=30'd781608573;
array[274]=30'd856066696;
array[275]=30'd856066696;
array[276]=30'd824623759;
array[277]=30'd814111379;
array[278]=30'd824623759;
array[279]=30'd824623759;
array[280]=30'd856066696;
array[281]=30'd856066696;
array[282]=30'd856066696;
array[283]=30'd856066696;
array[284]=30'd856066696;
array[285]=30'd879168118;
array[286]=30'd898043496;
array[287]=30'd959928886;
array[288]=30'd856066696;
array[289]=30'd856066696;
array[290]=30'd856066696;
array[291]=30'd856066696;
array[292]=30'd856066696;
array[293]=30'd856066696;
array[294]=30'd841408084;
array[295]=30'd739680847;
array[296]=30'd428280389;
array[297]=30'd439849468;
array[298]=30'd709306968;
array[299]=30'd856066696;
array[300]=30'd856066696;
array[301]=30'd856066696;
array[302]=30'd856066696;
array[303]=30'd856066696;
array[304]=30'd856066696;
array[305]=30'd856066696;
array[306]=30'd856066696;
array[307]=30'd856066696;
array[308]=30'd856066696;
array[309]=30'd856066696;
array[310]=30'd856066696;
array[311]=30'd856066696;
array[312]=30'd856066696;
array[313]=30'd856066696;
array[314]=30'd856066696;
array[315]=30'd856066696;
array[316]=30'd856066696;
array[317]=30'd856066696;
array[318]=30'd856066696;
array[319]=30'd856066696;
array[320]=30'd856066696;
array[321]=30'd856066696;
array[322]=30'd856066696;
array[323]=30'd856066696;
array[324]=30'd856066696;
array[325]=30'd856066696;
array[326]=30'd856066696;
array[327]=30'd856066696;
array[328]=30'd856066696;
array[329]=30'd856066696;
array[330]=30'd653676161;
array[331]=30'd467006094;
array[332]=30'd551919254;
array[333]=30'd559255224;
array[334]=30'd559255224;
array[335]=30'd608527024;
array[336]=30'd516257448;
array[337]=30'd646262454;
array[338]=30'd646262454;
array[339]=30'd516257448;
array[340]=30'd551919254;
array[341]=30'd633661142;
array[342]=30'd633661142;
array[343]=30'd582343294;
array[344]=30'd938933826;
array[345]=30'd841408084;
array[346]=30'd559303250;
array[347]=30'd634745492;
array[348]=30'd581260986;
array[349]=30'd633661142;
array[350]=30'd650433234;
array[351]=30'd608527024;
array[352]=30'd559255224;
array[353]=30'd633661142;
array[354]=30'd633661142;
array[355]=30'd633661142;
array[356]=30'd650433234;
array[357]=30'd633661142;
array[358]=30'd581260986;
array[359]=30'd310773397;
array[360]=30'd559255224;
array[361]=30'd633661142;
array[362]=30'd633661142;
array[363]=30'd633661142;
array[364]=30'd646262454;
array[365]=30'd559255224;
array[366]=30'd633661142;
array[367]=30'd646262454;
array[368]=30'd559255224;
array[369]=30'd781608573;
array[370]=30'd856066696;
array[371]=30'd824623759;
array[372]=30'd856066696;
array[373]=30'd824623759;
array[374]=30'd824623759;
array[375]=30'd856066696;
array[376]=30'd856066696;
array[377]=30'd856066696;
array[378]=30'd856066696;
array[379]=30'd856066696;
array[380]=30'd898043496;
array[381]=30'd959928886;
array[382]=30'd1000848926;
array[383]=30'd921177592;
array[384]=30'd856066696;
array[385]=30'd856066696;
array[386]=30'd856066696;
array[387]=30'd856066696;
array[388]=30'd824623759;
array[389]=30'd794241637;
array[390]=30'd597116464;
array[391]=30'd401043987;
array[392]=30'd456626661;
array[393]=30'd477594065;
array[394]=30'd439849468;
array[395]=30'd795279924;
array[396]=30'd856066696;
array[397]=30'd856066696;
array[398]=30'd856066696;
array[399]=30'd856066696;
array[400]=30'd856066696;
array[401]=30'd856066696;
array[402]=30'd856066696;
array[403]=30'd856066696;
array[404]=30'd856066696;
array[405]=30'd856066696;
array[406]=30'd856066696;
array[407]=30'd856066696;
array[408]=30'd856066696;
array[409]=30'd856066696;
array[410]=30'd856066696;
array[411]=30'd856066696;
array[412]=30'd856066696;
array[413]=30'd856066696;
array[414]=30'd856066696;
array[415]=30'd856066696;
array[416]=30'd856066696;
array[417]=30'd856066696;
array[418]=30'd856066696;
array[419]=30'd856066696;
array[420]=30'd856066696;
array[421]=30'd856066696;
array[422]=30'd856066696;
array[423]=30'd856066696;
array[424]=30'd856066696;
array[425]=30'd814111379;
array[426]=30'd496374434;
array[427]=30'd467006094;
array[428]=30'd634745492;
array[429]=30'd496374434;
array[430]=30'd608527024;
array[431]=30'd559255224;
array[432]=30'd559255224;
array[433]=30'd646262454;
array[434]=30'd646262454;
array[435]=30'd496374434;
array[436]=30'd559255224;
array[437]=30'd646262454;
array[438]=30'd608527024;
array[439]=30'd739680847;
array[440]=30'd938933826;
array[441]=30'd884420162;
array[442]=30'd527847013;
array[443]=30'd634745492;
array[444]=30'd444952244;
array[445]=30'd608527024;
array[446]=30'd646262454;
array[447]=30'd646262454;
array[448]=30'd427157133;
array[449]=30'd646262454;
array[450]=30'd633661142;
array[451]=30'd633661142;
array[452]=30'd633661142;
array[453]=30'd608527024;
array[454]=30'd608527024;
array[455]=30'd310773397;
array[456]=30'd522581659;
array[457]=30'd633661142;
array[458]=30'd633661142;
array[459]=30'd633661142;
array[460]=30'd650433234;
array[461]=30'd516257448;
array[462]=30'd646262454;
array[463]=30'd646262454;
array[464]=30'd608527024;
array[465]=30'd686214797;
array[466]=30'd856066696;
array[467]=30'd856066696;
array[468]=30'd824623759;
array[469]=30'd814111379;
array[470]=30'd856066696;
array[471]=30'd856066696;
array[472]=30'd856066696;
array[473]=30'd856066696;
array[474]=30'd856066696;
array[475]=30'd856066696;
array[476]=30'd884420162;
array[477]=30'd855119431;
array[478]=30'd785935846;
array[479]=30'd758671804;
array[480]=30'd856066696;
array[481]=30'd856066696;
array[482]=30'd856066696;
array[483]=30'd856066696;
array[484]=30'd794241637;
array[485]=30'd506974798;
array[486]=30'd341289472;
array[487]=30'd439849468;
array[488]=30'd396870070;
array[489]=30'd472369584;
array[490]=30'd425179585;
array[491]=30'd617030138;
array[492]=30'd841408084;
array[493]=30'd879168118;
array[494]=30'd879168118;
array[495]=30'd841408084;
array[496]=30'd841408084;
array[497]=30'd841408084;
array[498]=30'd841408084;
array[499]=30'd856066696;
array[500]=30'd879168118;
array[501]=30'd841408084;
array[502]=30'd841408084;
array[503]=30'd856066696;
array[504]=30'd856066696;
array[505]=30'd856066696;
array[506]=30'd856066696;
array[507]=30'd856066696;
array[508]=30'd856066696;
array[509]=30'd856066696;
array[510]=30'd856066696;
array[511]=30'd856066696;
array[512]=30'd856066696;
array[513]=30'd856066696;
array[514]=30'd856066696;
array[515]=30'd856066696;
array[516]=30'd856066696;
array[517]=30'd856066696;
array[518]=30'd856066696;
array[519]=30'd856066696;
array[520]=30'd824623759;
array[521]=30'd729186945;
array[522]=30'd483822211;
array[523]=30'd467006094;
array[524]=30'd646262454;
array[525]=30'd444952244;
array[526]=30'd646262454;
array[527]=30'd516257448;
array[528]=30'd608527024;
array[529]=30'd646262454;
array[530]=30'd559255224;
array[531]=30'd605405812;
array[532]=30'd582343294;
array[533]=30'd646262454;
array[534]=30'd551919254;
array[535]=30'd884420162;
array[536]=30'd938933826;
array[537]=30'd884420162;
array[538]=30'd496412259;
array[539]=30'd605405812;
array[540]=30'd605405812;
array[541]=30'd558250630;
array[542]=30'd646262454;
array[543]=30'd646262454;
array[544]=30'd496374434;
array[545]=30'd551919254;
array[546]=30'd646262454;
array[547]=30'd633661142;
array[548]=30'd633661142;
array[549]=30'd516257448;
array[550]=30'd608527024;
array[551]=30'd340142721;
array[552]=30'd467006094;
array[553]=30'd646262454;
array[554]=30'd633661142;
array[555]=30'd633661142;
array[556]=30'd633661142;
array[557]=30'd608527024;
array[558]=30'd547692230;
array[559]=30'd633661142;
array[560]=30'd646262454;
array[561]=30'd613805729;
array[562]=30'd856066696;
array[563]=30'd856066696;
array[564]=30'd856066696;
array[565]=30'd856066696;
array[566]=30'd856066696;
array[567]=30'd856066696;
array[568]=30'd856066696;
array[569]=30'd856066696;
array[570]=30'd856066696;
array[571]=30'd856066696;
array[572]=30'd879168118;
array[573]=30'd810005031;
array[574]=30'd810005031;
array[575]=30'd821544417;
array[576]=30'd856066696;
array[577]=30'd856066696;
array[578]=30'd856066696;
array[579]=30'd856066696;
array[580]=30'd744990312;
array[581]=30'd401043987;
array[582]=30'd456626661;
array[583]=30'd343392696;
array[584]=30'd425179585;
array[585]=30'd472369584;
array[586]=30'd472369584;
array[587]=30'd456626661;
array[588]=30'd843548160;
array[589]=30'd903304711;
array[590]=30'd860309028;
array[591]=30'd843548160;
array[592]=30'd843548160;
array[593]=30'd843548160;
array[594]=30'd810005031;
array[595]=30'd597116464;
array[596]=30'd597116464;
array[597]=30'd843548160;
array[598]=30'd843548160;
array[599]=30'd860309028;
array[600]=30'd856066696;
array[601]=30'd856066696;
array[602]=30'd856066696;
array[603]=30'd856066696;
array[604]=30'd856066696;
array[605]=30'd856066696;
array[606]=30'd856066696;
array[607]=30'd856066696;
array[608]=30'd856066696;
array[609]=30'd856066696;
array[610]=30'd856066696;
array[611]=30'd856066696;
array[612]=30'd856066696;
array[613]=30'd856066696;
array[614]=30'd856066696;
array[615]=30'd824623759;
array[616]=30'd824623759;
array[617]=30'd582343294;
array[618]=30'd558250630;
array[619]=30'd522581659;
array[620]=30'd646262454;
array[621]=30'd485848753;
array[622]=30'd646262454;
array[623]=30'd427157133;
array[624]=30'd608527024;
array[625]=30'd608527024;
array[626]=30'd558250630;
array[627]=30'd709306968;
array[628]=30'd605405812;
array[629]=30'd608527024;
array[630]=30'd624350812;
array[631]=30'd938933826;
array[632]=30'd959928886;
array[633]=30'd916921900;
array[634]=30'd537304625;
array[635]=30'd605405812;
array[636]=30'd756500033;
array[637]=30'd527847013;
array[638]=30'd634745492;
array[639]=30'd646262454;
array[640]=30'd653676161;
array[641]=30'd592910950;
array[642]=30'd634745492;
array[643]=30'd646262454;
array[644]=30'd646262454;
array[645]=30'd444952244;
array[646]=30'd559255224;
array[647]=30'd387329638;
array[648]=30'd408333955;
array[649]=30'd646262454;
array[650]=30'd633661142;
array[651]=30'd633661142;
array[652]=30'd633661142;
array[653]=30'd633661142;
array[654]=30'd516257448;
array[655]=30'd633661142;
array[656]=30'd646262454;
array[657]=30'd551919254;
array[658]=30'd856066696;
array[659]=30'd856066696;
array[660]=30'd824623759;
array[661]=30'd824623759;
array[662]=30'd856066696;
array[663]=30'd856066696;
array[664]=30'd856066696;
array[665]=30'd856066696;
array[666]=30'd856066696;
array[667]=30'd856066696;
array[668]=30'd856066696;
array[669]=30'd879168118;
array[670]=30'd841408084;
array[671]=30'd841408084;
array[672]=30'd856066696;
array[673]=30'd856066696;
array[674]=30'd856066696;
array[675]=30'd856066696;
array[676]=30'd841408084;
array[677]=30'd458750516;
array[678]=30'd484957641;
array[679]=30'd396870070;
array[680]=30'd425179585;
array[681]=30'd472369584;
array[682]=30'd472369584;
array[683]=30'd472369584;
array[684]=30'd541585861;
array[685]=30'd774396326;
array[686]=30'd758671804;
array[687]=30'd740853147;
array[688]=30'd774396326;
array[689]=30'd758671804;
array[690]=30'd740803022;
array[691]=30'd396870070;
array[692]=30'd425179585;
array[693]=30'd621275606;
array[694]=30'd798493124;
array[695]=30'd843548160;
array[696]=30'd841408084;
array[697]=30'd856066696;
array[698]=30'd856066696;
array[699]=30'd856066696;
array[700]=30'd856066696;
array[701]=30'd856066696;
array[702]=30'd856066696;
array[703]=30'd856066696;
array[704]=30'd856066696;
array[705]=30'd856066696;
array[706]=30'd856066696;
array[707]=30'd856066696;
array[708]=30'd856066696;
array[709]=30'd856066696;
array[710]=30'd856066696;
array[711]=30'd856066696;
array[712]=30'd795279924;
array[713]=30'd448143984;
array[714]=30'd558250630;
array[715]=30'd551919254;
array[716]=30'd608527024;
array[717]=30'd452327079;
array[718]=30'd608527024;
array[719]=30'd331722417;
array[720]=30'd634745492;
array[721]=30'd608527024;
array[722]=30'd624350812;
array[723]=30'd795279924;
array[724]=30'd582343294;
array[725]=30'd634745492;
array[726]=30'd739680847;
array[727]=30'd959928886;
array[728]=30'd938933826;
array[729]=30'd938933826;
array[730]=30'd624350812;
array[731]=30'd592910950;
array[732]=30'd815194717;
array[733]=30'd756500033;
array[734]=30'd582343294;
array[735]=30'd646262454;
array[736]=30'd558250630;
array[737]=30'd756500033;
array[738]=30'd582343294;
array[739]=30'd608527024;
array[740]=30'd646262454;
array[741]=30'd551919254;
array[742]=30'd522581659;
array[743]=30'd448143984;
array[744]=30'd387329638;
array[745]=30'd634745492;
array[746]=30'd646262454;
array[747]=30'd633661142;
array[748]=30'd633661142;
array[749]=30'd633661142;
array[750]=30'd516257448;
array[751]=30'd633661142;
array[752]=30'd646262454;
array[753]=30'd516257448;
array[754]=30'd814111379;
array[755]=30'd856066696;
array[756]=30'd856066696;
array[757]=30'd824623759;
array[758]=30'd856066696;
array[759]=30'd856066696;
array[760]=30'd856066696;
array[761]=30'd856066696;
array[762]=30'd856066696;
array[763]=30'd856066696;
array[764]=30'd856066696;
array[765]=30'd856066696;
array[766]=30'd856066696;
array[767]=30'd879168118;
array[768]=30'd856066696;
array[769]=30'd856066696;
array[770]=30'd856066696;
array[771]=30'd856066696;
array[772]=30'd879168118;
array[773]=30'd725091917;
array[774]=30'd383250907;
array[775]=30'd472369584;
array[776]=30'd396870070;
array[777]=30'd491240873;
array[778]=30'd472369584;
array[779]=30'd472369584;
array[780]=30'd425179585;
array[781]=30'd816348600;
array[782]=30'd911766951;
array[783]=30'd790145435;
array[784]=30'd850952611;
array[785]=30'd911766951;
array[786]=30'd674763200;
array[787]=30'd425179585;
array[788]=30'd472369584;
array[789]=30'd484957641;
array[790]=30'd798493124;
array[791]=30'd821544417;
array[792]=30'd860309028;
array[793]=30'd824623759;
array[794]=30'd856066696;
array[795]=30'd856066696;
array[796]=30'd856066696;
array[797]=30'd856066696;
array[798]=30'd856066696;
array[799]=30'd856066696;
array[800]=30'd856066696;
array[801]=30'd856066696;
array[802]=30'd856066696;
array[803]=30'd856066696;
array[804]=30'd856066696;
array[805]=30'd856066696;
array[806]=30'd856066696;
array[807]=30'd879168118;
array[808]=30'd815194717;
array[809]=30'd485876339;
array[810]=30'd582343294;
array[811]=30'd551919254;
array[812]=30'd608527024;
array[813]=30'd362130088;
array[814]=30'd551919254;
array[815]=30'd434534016;
array[816]=30'd605405812;
array[817]=30'd559255224;
array[818]=30'd739680847;
array[819]=30'd795279924;
array[820]=30'd527847013;
array[821]=30'd582343294;
array[822]=30'd841408084;
array[823]=30'd959928886;
array[824]=30'd938933826;
array[825]=30'd938933826;
array[826]=30'd795279924;
array[827]=30'd527847013;
array[828]=30'd795279924;
array[829]=30'd916921900;
array[830]=30'd527847013;
array[831]=30'd634745492;
array[832]=30'd483822211;
array[833]=30'd884420162;
array[834]=30'd527847013;
array[835]=30'd634745492;
array[836]=30'd608527024;
array[837]=30'd582343294;
array[838]=30'd527847013;
array[839]=30'd592910950;
array[840]=30'd459725411;
array[841]=30'd634745492;
array[842]=30'd646262454;
array[843]=30'd633661142;
array[844]=30'd633661142;
array[845]=30'd633661142;
array[846]=30'd559255224;
array[847]=30'd646262454;
array[848]=30'd633661142;
array[849]=30'd551919254;
array[850]=30'd781608573;
array[851]=30'd856066696;
array[852]=30'd856066696;
array[853]=30'd824623759;
array[854]=30'd856066696;
array[855]=30'd856066696;
array[856]=30'd856066696;
array[857]=30'd856066696;
array[858]=30'd856066696;
array[859]=30'd856066696;
array[860]=30'd856066696;
array[861]=30'd856066696;
array[862]=30'd856066696;
array[863]=30'd879168118;
array[864]=30'd856066696;
array[865]=30'd856066696;
array[866]=30'd856066696;
array[867]=30'd856066696;
array[868]=30'd856066696;
array[869]=30'd842499661;
array[870]=30'd528973367;
array[871]=30'd456626661;
array[872]=30'd396870070;
array[873]=30'd472369584;
array[874]=30'd491240873;
array[875]=30'd491240873;
array[876]=30'd472369584;
array[877]=30'd642253230;
array[878]=30'd790145435;
array[879]=30'd740853147;
array[880]=30'd774396326;
array[881]=30'd945316283;
array[882]=30'd592970169;
array[883]=30'd472369584;
array[884]=30'd472369584;
array[885]=30'd343392696;
array[886]=30'd642253230;
array[887]=30'd758671804;
array[888]=30'd843548160;
array[889]=30'd841408084;
array[890]=30'd856066696;
array[891]=30'd856066696;
array[892]=30'd856066696;
array[893]=30'd856066696;
array[894]=30'd856066696;
array[895]=30'd856066696;
array[896]=30'd856066696;
array[897]=30'd856066696;
array[898]=30'd856066696;
array[899]=30'd856066696;
array[900]=30'd856066696;
array[901]=30'd856066696;
array[902]=30'd856066696;
array[903]=30'd879168118;
array[904]=30'd795279924;
array[905]=30'd559303250;
array[906]=30'd605405812;
array[907]=30'd522581659;
array[908]=30'd613805729;
array[909]=30'd340142721;
array[910]=30'd527847013;
array[911]=30'd624350812;
array[912]=30'd582343294;
array[913]=30'd527847013;
array[914]=30'd665233987;
array[915]=30'd795279924;
array[916]=30'd512140869;
array[917]=30'd496412259;
array[918]=30'd795279924;
array[919]=30'd959928886;
array[920]=30'd959928886;
array[921]=30'd959928886;
array[922]=30'd884420162;
array[923]=30'd512140869;
array[924]=30'd668430907;
array[925]=30'd694642226;
array[926]=30'd712431145;
array[927]=30'd558250630;
array[928]=30'd496412259;
array[929]=30'd665233987;
array[930]=30'd624350812;
array[931]=30'd582343294;
array[932]=30'd634745492;
array[933]=30'd592910950;
array[934]=30'd566698607;
array[935]=30'd597116464;
array[936]=30'd665233987;
array[937]=30'd625322602;
array[938]=30'd646262454;
array[939]=30'd608527024;
array[940]=30'd646262454;
array[941]=30'd633661142;
array[942]=30'd547692230;
array[943]=30'd581260986;
array[944]=30'd646262454;
array[945]=30'd559255224;
array[946]=30'd781608573;
array[947]=30'd856066696;
array[948]=30'd856066696;
array[949]=30'd856066696;
array[950]=30'd856066696;
array[951]=30'd856066696;
array[952]=30'd856066696;
array[953]=30'd856066696;
array[954]=30'd856066696;
array[955]=30'd856066696;
array[956]=30'd856066696;
array[957]=30'd856066696;
array[958]=30'd856066696;
array[959]=30'd879168118;
array[960]=30'd856066696;
array[961]=30'd856066696;
array[962]=30'd856066696;
array[963]=30'd856066696;
array[964]=30'd856066696;
array[965]=30'd879168118;
array[966]=30'd744990312;
array[967]=30'd426248712;
array[968]=30'd463997419;
array[969]=30'd425179585;
array[970]=30'd472369584;
array[971]=30'd491240873;
array[972]=30'd472369584;
array[973]=30'd425179585;
array[974]=30'd758671804;
array[975]=30'd816348600;
array[976]=30'd774396326;
array[977]=30'd945316283;
array[978]=30'd425179585;
array[979]=30'd472369584;
array[980]=30'd472369584;
array[981]=30'd396870070;
array[982]=30'd425179585;
array[983]=30'd674763200;
array[984]=30'd843548160;
array[985]=30'd841408084;
array[986]=30'd856066696;
array[987]=30'd856066696;
array[988]=30'd856066696;
array[989]=30'd856066696;
array[990]=30'd856066696;
array[991]=30'd856066696;
array[992]=30'd856066696;
array[993]=30'd856066696;
array[994]=30'd856066696;
array[995]=30'd856066696;
array[996]=30'd856066696;
array[997]=30'd856066696;
array[998]=30'd856066696;
array[999]=30'd879168118;
array[1000]=30'd683036269;
array[1001]=30'd605405812;
array[1002]=30'd613805729;
array[1003]=30'd496374434;
array[1004]=30'd559255224;
array[1005]=30'd483822211;
array[1006]=30'd496412259;
array[1007]=30'd795279924;
array[1008]=30'd459725411;
array[1009]=30'd559303250;
array[1010]=30'd938933826;
array[1011]=30'd938933826;
array[1012]=30'd694642226;
array[1013]=30'd496412259;
array[1014]=30'd938933826;
array[1015]=30'd979842606;
array[1016]=30'd959928886;
array[1017]=30'd959928886;
array[1018]=30'd938933826;
array[1019]=30'd756500033;
array[1020]=30'd694642226;
array[1021]=30'd959928886;
array[1022]=30'd938933826;
array[1023]=30'd624350812;
array[1024]=30'd527847013;
array[1025]=30'd916921900;
array[1026]=30'd860309028;
array[1027]=30'd527847013;
array[1028]=30'd605405812;
array[1029]=30'd668430907;
array[1030]=30'd668430907;
array[1031]=30'd668430907;
array[1032]=30'd756500033;
array[1033]=30'd582343294;
array[1034]=30'd608527024;
array[1035]=30'd581260986;
array[1036]=30'd608527024;
array[1037]=30'd633661142;
array[1038]=30'd581260986;
array[1039]=30'd559255224;
array[1040]=30'd633661142;
array[1041]=30'd581260986;
array[1042]=30'd729186945;
array[1043]=30'd856066696;
array[1044]=30'd856066696;
array[1045]=30'd856066696;
array[1046]=30'd856066696;
array[1047]=30'd856066696;
array[1048]=30'd856066696;
array[1049]=30'd856066696;
array[1050]=30'd856066696;
array[1051]=30'd856066696;
array[1052]=30'd856066696;
array[1053]=30'd856066696;
array[1054]=30'd856066696;
array[1055]=30'd856066696;
array[1056]=30'd856066696;
array[1057]=30'd856066696;
array[1058]=30'd856066696;
array[1059]=30'd856066696;
array[1060]=30'd856066696;
array[1061]=30'd879168118;
array[1062]=30'd879168118;
array[1063]=30'd612873765;
array[1064]=30'd426248712;
array[1065]=30'd472369584;
array[1066]=30'd491240873;
array[1067]=30'd491240873;
array[1068]=30'd491240873;
array[1069]=30'd472369584;
array[1070]=30'd621275606;
array[1071]=30'd945316283;
array[1072]=30'd871910847;
array[1073]=30'd798493124;
array[1074]=30'd396870070;
array[1075]=30'd472369584;
array[1076]=30'd425179585;
array[1077]=30'd425179585;
array[1078]=30'd425179585;
array[1079]=30'd674763200;
array[1080]=30'd843548160;
array[1081]=30'd841408084;
array[1082]=30'd856066696;
array[1083]=30'd856066696;
array[1084]=30'd856066696;
array[1085]=30'd856066696;
array[1086]=30'd856066696;
array[1087]=30'd856066696;
array[1088]=30'd856066696;
array[1089]=30'd856066696;
array[1090]=30'd856066696;
array[1091]=30'd856066696;
array[1092]=30'd856066696;
array[1093]=30'd856066696;
array[1094]=30'd856066696;
array[1095]=30'd856066696;
array[1096]=30'd624350812;
array[1097]=30'd634745492;
array[1098]=30'd608527024;
array[1099]=30'd444952244;
array[1100]=30'd559255224;
array[1101]=30'd709306968;
array[1102]=30'd428280389;
array[1103]=30'd712431145;
array[1104]=30'd582384191;
array[1105]=30'd548890196;
array[1106]=30'd959928886;
array[1107]=30'd959928886;
array[1108]=30'd884420162;
array[1109]=30'd571952708;
array[1110]=30'd959928886;
array[1111]=30'd959928886;
array[1112]=30'd959928886;
array[1113]=30'd959928886;
array[1114]=30'd959928886;
array[1115]=30'd916921900;
array[1116]=30'd795279924;
array[1117]=30'd979842606;
array[1118]=30'd959928886;
array[1119]=30'd884420162;
array[1120]=30'd537304625;
array[1121]=30'd916921900;
array[1122]=30'd959928886;
array[1123]=30'd739680847;
array[1124]=30'd459725411;
array[1125]=30'd756500033;
array[1126]=30'd725052963;
array[1127]=30'd756500033;
array[1128]=30'd756500033;
array[1129]=30'd512140869;
array[1130]=30'd634745492;
array[1131]=30'd559255224;
array[1132]=30'd608527024;
array[1133]=30'd646262454;
array[1134]=30'd646262454;
array[1135]=30'd559255224;
array[1136]=30'd633661142;
array[1137]=30'd608527024;
array[1138]=30'd729186945;
array[1139]=30'd856066696;
array[1140]=30'd856066696;
array[1141]=30'd856066696;
array[1142]=30'd856066696;
array[1143]=30'd856066696;
array[1144]=30'd856066696;
array[1145]=30'd856066696;
array[1146]=30'd856066696;
array[1147]=30'd856066696;
array[1148]=30'd856066696;
array[1149]=30'd856066696;
array[1150]=30'd856066696;
array[1151]=30'd856066696;
array[1152]=30'd856066696;
array[1153]=30'd856066696;
array[1154]=30'd856066696;
array[1155]=30'd856066696;
array[1156]=30'd856066696;
array[1157]=30'd879168118;
array[1158]=30'd879168118;
array[1159]=30'd842499661;
array[1160]=30'd458750516;
array[1161]=30'd477594065;
array[1162]=30'd472369584;
array[1163]=30'd491240873;
array[1164]=30'd491240873;
array[1165]=30'd472369584;
array[1166]=30'd472369584;
array[1167]=30'd945316283;
array[1168]=30'd816348600;
array[1169]=30'd541585861;
array[1170]=30'd425179585;
array[1171]=30'd472369584;
array[1172]=30'd396870070;
array[1173]=30'd472369584;
array[1174]=30'd396870070;
array[1175]=30'd740803022;
array[1176]=30'd860309028;
array[1177]=30'd856066696;
array[1178]=30'd856066696;
array[1179]=30'd856066696;
array[1180]=30'd856066696;
array[1181]=30'd856066696;
array[1182]=30'd856066696;
array[1183]=30'd856066696;
array[1184]=30'd856066696;
array[1185]=30'd856066696;
array[1186]=30'd856066696;
array[1187]=30'd856066696;
array[1188]=30'd856066696;
array[1189]=30'd856066696;
array[1190]=30'd856066696;
array[1191]=30'd856066696;
array[1192]=30'd592910950;
array[1193]=30'd634745492;
array[1194]=30'd646262454;
array[1195]=30'd516257448;
array[1196]=30'd522581659;
array[1197]=30'd709306968;
array[1198]=30'd428280389;
array[1199]=30'd916921900;
array[1200]=30'd884420162;
array[1201]=30'd571952708;
array[1202]=30'd959928886;
array[1203]=30'd959928886;
array[1204]=30'd959928886;
array[1205]=30'd916921900;
array[1206]=30'd959928886;
array[1207]=30'd959928886;
array[1208]=30'd959928886;
array[1209]=30'd959928886;
array[1210]=30'd959928886;
array[1211]=30'd959928886;
array[1212]=30'd959928886;
array[1213]=30'd959928886;
array[1214]=30'd959928886;
array[1215]=30'd959928886;
array[1216]=30'd884420162;
array[1217]=30'd938933826;
array[1218]=30'd959928886;
array[1219]=30'd884420162;
array[1220]=30'd512140869;
array[1221]=30'd860309028;
array[1222]=30'd597116464;
array[1223]=30'd810005031;
array[1224]=30'd439849468;
array[1225]=30'd475488805;
array[1226]=30'd448143984;
array[1227]=30'd522581659;
array[1228]=30'd608527024;
array[1229]=30'd633661142;
array[1230]=30'd646262454;
array[1231]=30'd547692230;
array[1232]=30'd650433234;
array[1233]=30'd581260986;
array[1234]=30'd729186945;
array[1235]=30'd856066696;
array[1236]=30'd856066696;
array[1237]=30'd856066696;
array[1238]=30'd856066696;
array[1239]=30'd856066696;
array[1240]=30'd856066696;
array[1241]=30'd856066696;
array[1242]=30'd856066696;
array[1243]=30'd856066696;
array[1244]=30'd856066696;
array[1245]=30'd856066696;
array[1246]=30'd856066696;
array[1247]=30'd856066696;
array[1248]=30'd856066696;
array[1249]=30'd856066696;
array[1250]=30'd856066696;
array[1251]=30'd856066696;
array[1252]=30'd879168118;
array[1253]=30'd879168118;
array[1254]=30'd879168118;
array[1255]=30'd879168118;
array[1256]=30'd709306968;
array[1257]=30'd439849468;
array[1258]=30'd472369584;
array[1259]=30'd472369584;
array[1260]=30'd491240873;
array[1261]=30'd491240873;
array[1262]=30'd425179585;
array[1263]=30'd621275606;
array[1264]=30'd740853147;
array[1265]=30'd396870070;
array[1266]=30'd472369584;
array[1267]=30'd472369584;
array[1268]=30'd425179585;
array[1269]=30'd472369584;
array[1270]=30'd396870070;
array[1271]=30'd843548160;
array[1272]=30'd841408084;
array[1273]=30'd856066696;
array[1274]=30'd856066696;
array[1275]=30'd856066696;
array[1276]=30'd856066696;
array[1277]=30'd856066696;
array[1278]=30'd856066696;
array[1279]=30'd856066696;
array[1280]=30'd856066696;
array[1281]=30'd856066696;
array[1282]=30'd856066696;
array[1283]=30'd856066696;
array[1284]=30'd856066696;
array[1285]=30'd856066696;
array[1286]=30'd856066696;
array[1287]=30'd856066696;
array[1288]=30'd558250630;
array[1289]=30'd634745492;
array[1290]=30'd646262454;
array[1291]=30'd608527024;
array[1292]=30'd427157133;
array[1293]=30'd756500033;
array[1294]=30'd860309028;
array[1295]=30'd959928886;
array[1296]=30'd959928886;
array[1297]=30'd884420162;
array[1298]=30'd959928886;
array[1299]=30'd959928886;
array[1300]=30'd959928886;
array[1301]=30'd959928886;
array[1302]=30'd959928886;
array[1303]=30'd959928886;
array[1304]=30'd959928886;
array[1305]=30'd979842606;
array[1306]=30'd959928886;
array[1307]=30'd959928886;
array[1308]=30'd979842606;
array[1309]=30'd979842606;
array[1310]=30'd959928886;
array[1311]=30'd959928886;
array[1312]=30'd959928886;
array[1313]=30'd959928886;
array[1314]=30'd959928886;
array[1315]=30'd959928886;
array[1316]=30'd916921900;
array[1317]=30'd959928886;
array[1318]=30'd860309028;
array[1319]=30'd810005031;
array[1320]=30'd649571855;
array[1321]=30'd821544417;
array[1322]=30'd462859830;
array[1323]=30'd485876339;
array[1324]=30'd634745492;
array[1325]=30'd646262454;
array[1326]=30'd646262454;
array[1327]=30'd547692230;
array[1328]=30'd650433234;
array[1329]=30'd581260986;
array[1330]=30'd781608573;
array[1331]=30'd856066696;
array[1332]=30'd856066696;
array[1333]=30'd856066696;
array[1334]=30'd856066696;
array[1335]=30'd856066696;
array[1336]=30'd856066696;
array[1337]=30'd856066696;
array[1338]=30'd856066696;
array[1339]=30'd856066696;
array[1340]=30'd856066696;
array[1341]=30'd856066696;
array[1342]=30'd856066696;
array[1343]=30'd856066696;
array[1344]=30'd856066696;
array[1345]=30'd856066696;
array[1346]=30'd856066696;
array[1347]=30'd856066696;
array[1348]=30'd856066696;
array[1349]=30'd856066696;
array[1350]=30'd879168118;
array[1351]=30'd879168118;
array[1352]=30'd842499661;
array[1353]=30'd555187752;
array[1354]=30'd463997419;
array[1355]=30'd491240873;
array[1356]=30'd491240873;
array[1357]=30'd491240873;
array[1358]=30'd472369584;
array[1359]=30'd425179585;
array[1360]=30'd758671804;
array[1361]=30'd396870070;
array[1362]=30'd472369584;
array[1363]=30'd472369584;
array[1364]=30'd472369584;
array[1365]=30'd425179585;
array[1366]=30'd477594065;
array[1367]=30'd860309028;
array[1368]=30'd856066696;
array[1369]=30'd856066696;
array[1370]=30'd856066696;
array[1371]=30'd856066696;
array[1372]=30'd856066696;
array[1373]=30'd856066696;
array[1374]=30'd856066696;
array[1375]=30'd856066696;
array[1376]=30'd856066696;
array[1377]=30'd856066696;
array[1378]=30'd856066696;
array[1379]=30'd856066696;
array[1380]=30'd856066696;
array[1381]=30'd856066696;
array[1382]=30'd856066696;
array[1383]=30'd856066696;
array[1384]=30'd558250630;
array[1385]=30'd634745492;
array[1386]=30'd646262454;
array[1387]=30'd559255224;
array[1388]=30'd522581659;
array[1389]=30'd756500033;
array[1390]=30'd959928886;
array[1391]=30'd959928886;
array[1392]=30'd959928886;
array[1393]=30'd959928886;
array[1394]=30'd884420162;
array[1395]=30'd860309028;
array[1396]=30'd884420162;
array[1397]=30'd959928886;
array[1398]=30'd959928886;
array[1399]=30'd959928886;
array[1400]=30'd959928886;
array[1401]=30'd979842606;
array[1402]=30'd959928886;
array[1403]=30'd959928886;
array[1404]=30'd979842606;
array[1405]=30'd959928886;
array[1406]=30'd959928886;
array[1407]=30'd959928886;
array[1408]=30'd959928886;
array[1409]=30'd959928886;
array[1410]=30'd959928886;
array[1411]=30'd959928886;
array[1412]=30'd959928886;
array[1413]=30'd959928886;
array[1414]=30'd959928886;
array[1415]=30'd898098744;
array[1416]=30'd649571855;
array[1417]=30'd775423471;
array[1418]=30'd512140869;
array[1419]=30'd485876339;
array[1420]=30'd634745492;
array[1421]=30'd646262454;
array[1422]=30'd646262454;
array[1423]=30'd547692230;
array[1424]=30'd650433234;
array[1425]=30'd559255224;
array[1426]=30'd781608573;
array[1427]=30'd856066696;
array[1428]=30'd856066696;
array[1429]=30'd856066696;
array[1430]=30'd856066696;
array[1431]=30'd856066696;
array[1432]=30'd856066696;
array[1433]=30'd856066696;
array[1434]=30'd856066696;
array[1435]=30'd856066696;
array[1436]=30'd856066696;
array[1437]=30'd856066696;
array[1438]=30'd856066696;
array[1439]=30'd856066696;
array[1440]=30'd856066696;
array[1441]=30'd856066696;
array[1442]=30'd856066696;
array[1443]=30'd856066696;
array[1444]=30'd856066696;
array[1445]=30'd856066696;
array[1446]=30'd856066696;
array[1447]=30'd879168118;
array[1448]=30'd879168118;
array[1449]=30'd779606588;
array[1450]=30'd426248712;
array[1451]=30'd472369584;
array[1452]=30'd491240873;
array[1453]=30'd491240873;
array[1454]=30'd472369584;
array[1455]=30'd425179585;
array[1456]=30'd642253230;
array[1457]=30'd396870070;
array[1458]=30'd472369584;
array[1459]=30'd472369584;
array[1460]=30'd472369584;
array[1461]=30'd425179585;
array[1462]=30'd649571855;
array[1463]=30'd884420162;
array[1464]=30'd856066696;
array[1465]=30'd856066696;
array[1466]=30'd856066696;
array[1467]=30'd856066696;
array[1468]=30'd856066696;
array[1469]=30'd856066696;
array[1470]=30'd856066696;
array[1471]=30'd856066696;
array[1472]=30'd856066696;
array[1473]=30'd856066696;
array[1474]=30'd856066696;
array[1475]=30'd856066696;
array[1476]=30'd856066696;
array[1477]=30'd856066696;
array[1478]=30'd856066696;
array[1479]=30'd856066696;
array[1480]=30'd582343294;
array[1481]=30'd634745492;
array[1482]=30'd646262454;
array[1483]=30'd485848753;
array[1484]=30'd613805729;
array[1485]=30'd756500033;
array[1486]=30'd959928886;
array[1487]=30'd959928886;
array[1488]=30'd860309028;
array[1489]=30'd694642226;
array[1490]=30'd725052963;
array[1491]=30'd860309028;
array[1492]=30'd810005031;
array[1493]=30'd810005031;
array[1494]=30'd959928886;
array[1495]=30'd959928886;
array[1496]=30'd959928886;
array[1497]=30'd959928886;
array[1498]=30'd959928886;
array[1499]=30'd959928886;
array[1500]=30'd959928886;
array[1501]=30'd916921900;
array[1502]=30'd810005031;
array[1503]=30'd725052963;
array[1504]=30'd725052963;
array[1505]=30'd756500033;
array[1506]=30'd916921900;
array[1507]=30'd959928886;
array[1508]=30'd959928886;
array[1509]=30'd959928886;
array[1510]=30'd959928886;
array[1511]=30'd860309028;
array[1512]=30'd475488805;
array[1513]=30'd475488805;
array[1514]=30'd559303250;
array[1515]=30'd485876339;
array[1516]=30'd608527024;
array[1517]=30'd633661142;
array[1518]=30'd646262454;
array[1519]=30'd547692230;
array[1520]=30'd633661142;
array[1521]=30'd551919254;
array[1522]=30'd814111379;
array[1523]=30'd856066696;
array[1524]=30'd856066696;
array[1525]=30'd856066696;
array[1526]=30'd856066696;
array[1527]=30'd856066696;
array[1528]=30'd856066696;
array[1529]=30'd856066696;
array[1530]=30'd856066696;
array[1531]=30'd856066696;
array[1532]=30'd856066696;
array[1533]=30'd856066696;
array[1534]=30'd856066696;
array[1535]=30'd856066696;
array[1536]=30'd856066696;
array[1537]=30'd856066696;
array[1538]=30'd856066696;
array[1539]=30'd856066696;
array[1540]=30'd856066696;
array[1541]=30'd879168118;
array[1542]=30'd856066696;
array[1543]=30'd879168118;
array[1544]=30'd879168118;
array[1545]=30'd879168118;
array[1546]=30'd694642226;
array[1547]=30'd426248712;
array[1548]=30'd472369584;
array[1549]=30'd472369584;
array[1550]=30'd472369584;
array[1551]=30'd472369584;
array[1552]=30'd396870070;
array[1553]=30'd425179585;
array[1554]=30'd472369584;
array[1555]=30'd472369584;
array[1556]=30'd472369584;
array[1557]=30'd396870070;
array[1558]=30'd756500033;
array[1559]=30'd841408084;
array[1560]=30'd856066696;
array[1561]=30'd856066696;
array[1562]=30'd856066696;
array[1563]=30'd856066696;
array[1564]=30'd856066696;
array[1565]=30'd856066696;
array[1566]=30'd856066696;
array[1567]=30'd856066696;
array[1568]=30'd856066696;
array[1569]=30'd856066696;
array[1570]=30'd856066696;
array[1571]=30'd856066696;
array[1572]=30'd856066696;
array[1573]=30'd856066696;
array[1574]=30'd856066696;
array[1575]=30'd856066696;
array[1576]=30'd605405812;
array[1577]=30'd634745492;
array[1578]=30'd646262454;
array[1579]=30'd485848753;
array[1580]=30'd669371047;
array[1581]=30'd624350812;
array[1582]=30'd938933826;
array[1583]=30'd756500033;
array[1584]=30'd756500033;
array[1585]=30'd756500033;
array[1586]=30'd475488805;
array[1587]=30'd359106099;
array[1588]=30'd597116464;
array[1589]=30'd916921900;
array[1590]=30'd959928886;
array[1591]=30'd959928886;
array[1592]=30'd959928886;
array[1593]=30'd959928886;
array[1594]=30'd959928886;
array[1595]=30'd959928886;
array[1596]=30'd938933826;
array[1597]=30'd725052963;
array[1598]=30'd810005031;
array[1599]=30'd725052963;
array[1600]=30'd694642226;
array[1601]=30'd725052963;
array[1602]=30'd668430907;
array[1603]=30'd725052963;
array[1604]=30'd916921900;
array[1605]=30'd959928886;
array[1606]=30'd959928886;
array[1607]=30'd936883742;
array[1608]=30'd725052963;
array[1609]=30'd527847013;
array[1610]=30'd625322602;
array[1611]=30'd452327079;
array[1612]=30'd646262454;
array[1613]=30'd646262454;
array[1614]=30'd608527024;
array[1615]=30'd559255224;
array[1616]=30'd633661142;
array[1617]=30'd551919254;
array[1618]=30'd824623759;
array[1619]=30'd856066696;
array[1620]=30'd856066696;
array[1621]=30'd856066696;
array[1622]=30'd856066696;
array[1623]=30'd856066696;
array[1624]=30'd856066696;
array[1625]=30'd856066696;
array[1626]=30'd856066696;
array[1627]=30'd856066696;
array[1628]=30'd856066696;
array[1629]=30'd856066696;
array[1630]=30'd856066696;
array[1631]=30'd856066696;
array[1632]=30'd856066696;
array[1633]=30'd856066696;
array[1634]=30'd856066696;
array[1635]=30'd879168118;
array[1636]=30'd879168118;
array[1637]=30'd879168118;
array[1638]=30'd856066696;
array[1639]=30'd879168118;
array[1640]=30'd879168118;
array[1641]=30'd879168118;
array[1642]=30'd842499661;
array[1643]=30'd528973367;
array[1644]=30'd456626661;
array[1645]=30'd472369584;
array[1646]=30'd472369584;
array[1647]=30'd472369584;
array[1648]=30'd343392696;
array[1649]=30'd472369584;
array[1650]=30'd472369584;
array[1651]=30'd472369584;
array[1652]=30'd472369584;
array[1653]=30'd439849468;
array[1654]=30'd860309028;
array[1655]=30'd856066696;
array[1656]=30'd856066696;
array[1657]=30'd856066696;
array[1658]=30'd856066696;
array[1659]=30'd856066696;
array[1660]=30'd879168118;
array[1661]=30'd879168118;
array[1662]=30'd879168118;
array[1663]=30'd879168118;
array[1664]=30'd856066696;
array[1665]=30'd879168118;
array[1666]=30'd856066696;
array[1667]=30'd856066696;
array[1668]=30'd856066696;
array[1669]=30'd856066696;
array[1670]=30'd856066696;
array[1671]=30'd856066696;
array[1672]=30'd624350812;
array[1673]=30'd634745492;
array[1674]=30'd646262454;
array[1675]=30'd444952244;
array[1676]=30'd646262454;
array[1677]=30'd558250630;
array[1678]=30'd842499661;
array[1679]=30'd810005031;
array[1680]=30'd525850118;
array[1681]=30'd359106099;
array[1682]=30'd694642226;
array[1683]=30'd795279924;
array[1684]=30'd555187752;
array[1685]=30'd475488805;
array[1686]=30'd916921900;
array[1687]=30'd959928886;
array[1688]=30'd959928886;
array[1689]=30'd959928886;
array[1690]=30'd959928886;
array[1691]=30'd959928886;
array[1692]=30'd959928886;
array[1693]=30'd612873765;
array[1694]=30'd359106099;
array[1695]=30'd597116464;
array[1696]=30'd668430907;
array[1697]=30'd475488805;
array[1698]=30'd230137397;
array[1699]=30'd515315216;
array[1700]=30'd668430907;
array[1701]=30'd860309028;
array[1702]=30'd959928886;
array[1703]=30'd916921900;
array[1704]=30'd795279924;
array[1705]=30'd582343294;
array[1706]=30'd634745492;
array[1707]=30'd444952244;
array[1708]=30'd646262454;
array[1709]=30'd646262454;
array[1710]=30'd581260986;
array[1711]=30'd559255224;
array[1712]=30'd646262454;
array[1713]=30'd551919254;
array[1714]=30'd856066696;
array[1715]=30'd856066696;
array[1716]=30'd856066696;
array[1717]=30'd856066696;
array[1718]=30'd856066696;
array[1719]=30'd856066696;
array[1720]=30'd856066696;
array[1721]=30'd856066696;
array[1722]=30'd856066696;
array[1723]=30'd856066696;
array[1724]=30'd856066696;
array[1725]=30'd856066696;
array[1726]=30'd856066696;
array[1727]=30'd856066696;
array[1728]=30'd856066696;
array[1729]=30'd856066696;
array[1730]=30'd879168118;
array[1731]=30'd879168118;
array[1732]=30'd879168118;
array[1733]=30'd879168118;
array[1734]=30'd879168118;
array[1735]=30'd879168118;
array[1736]=30'd879168118;
array[1737]=30'd879168118;
array[1738]=30'd884420162;
array[1739]=30'd756500033;
array[1740]=30'd463997419;
array[1741]=30'd472369584;
array[1742]=30'd472369584;
array[1743]=30'd472369584;
array[1744]=30'd425179585;
array[1745]=30'd425179585;
array[1746]=30'd472369584;
array[1747]=30'd472369584;
array[1748]=30'd472369584;
array[1749]=30'd581396985;
array[1750]=30'd860309028;
array[1751]=30'd856066696;
array[1752]=30'd856066696;
array[1753]=30'd879168118;
array[1754]=30'd879168118;
array[1755]=30'd879168118;
array[1756]=30'd879168118;
array[1757]=30'd879168118;
array[1758]=30'd879168118;
array[1759]=30'd879168118;
array[1760]=30'd879168118;
array[1761]=30'd879168118;
array[1762]=30'd856066696;
array[1763]=30'd856066696;
array[1764]=30'd856066696;
array[1765]=30'd856066696;
array[1766]=30'd856066696;
array[1767]=30'd856066696;
array[1768]=30'd653676161;
array[1769]=30'd634745492;
array[1770]=30'd646262454;
array[1771]=30'd485848753;
array[1772]=30'd646262454;
array[1773]=30'd582343294;
array[1774]=30'd842499661;
array[1775]=30'd359106099;
array[1776]=30'd597116464;
array[1777]=30'd916921900;
array[1778]=30'd959928886;
array[1779]=30'd959928886;
array[1780]=30'd959928886;
array[1781]=30'd884420162;
array[1782]=30'd959928886;
array[1783]=30'd959928886;
array[1784]=30'd979842606;
array[1785]=30'd959928886;
array[1786]=30'd959928886;
array[1787]=30'd959928886;
array[1788]=30'd959928886;
array[1789]=30'd860309028;
array[1790]=30'd916921900;
array[1791]=30'd959928886;
array[1792]=30'd959928886;
array[1793]=30'd959928886;
array[1794]=30'd810005031;
array[1795]=30'd475488805;
array[1796]=30'd321370635;
array[1797]=30'd810005031;
array[1798]=30'd959928886;
array[1799]=30'd938933826;
array[1800]=30'd756500033;
array[1801]=30'd605405812;
array[1802]=30'd608527024;
array[1803]=30'd467006094;
array[1804]=30'd516257448;
array[1805]=30'd646262454;
array[1806]=30'd559255224;
array[1807]=30'd581260986;
array[1808]=30'd646262454;
array[1809]=30'd653676161;
array[1810]=30'd879168118;
array[1811]=30'd856066696;
array[1812]=30'd856066696;
array[1813]=30'd856066696;
array[1814]=30'd856066696;
array[1815]=30'd856066696;
array[1816]=30'd856066696;
array[1817]=30'd856066696;
array[1818]=30'd856066696;
array[1819]=30'd856066696;
array[1820]=30'd856066696;
array[1821]=30'd856066696;
array[1822]=30'd856066696;
array[1823]=30'd856066696;
array[1824]=30'd856066696;
array[1825]=30'd856066696;
array[1826]=30'd879168118;
array[1827]=30'd879168118;
array[1828]=30'd879168118;
array[1829]=30'd879168118;
array[1830]=30'd879168118;
array[1831]=30'd879168118;
array[1832]=30'd879168118;
array[1833]=30'd879168118;
array[1834]=30'd884420162;
array[1835]=30'd898098744;
array[1836]=30'd649571855;
array[1837]=30'd425179585;
array[1838]=30'd472369584;
array[1839]=30'd472369584;
array[1840]=30'd472369584;
array[1841]=30'd396870070;
array[1842]=30'd472369584;
array[1843]=30'd472369584;
array[1844]=30'd425179585;
array[1845]=30'd693598700;
array[1846]=30'd903304711;
array[1847]=30'd884420162;
array[1848]=30'd879168118;
array[1849]=30'd856066696;
array[1850]=30'd879168118;
array[1851]=30'd879168118;
array[1852]=30'd879168118;
array[1853]=30'd879168118;
array[1854]=30'd879168118;
array[1855]=30'd879168118;
array[1856]=30'd879168118;
array[1857]=30'd879168118;
array[1858]=30'd879168118;
array[1859]=30'd856066696;
array[1860]=30'd856066696;
array[1861]=30'd856066696;
array[1862]=30'd856066696;
array[1863]=30'd856066696;
array[1864]=30'd683036269;
array[1865]=30'd634745492;
array[1866]=30'd646262454;
array[1867]=30'd485848753;
array[1868]=30'd669371047;
array[1869]=30'd558250630;
array[1870]=30'd641178190;
array[1871]=30'd612873765;
array[1872]=30'd959928886;
array[1873]=30'd959928886;
array[1874]=30'd959928886;
array[1875]=30'd959928886;
array[1876]=30'd959928886;
array[1877]=30'd959928886;
array[1878]=30'd959928886;
array[1879]=30'd979842606;
array[1880]=30'd979842606;
array[1881]=30'd979842606;
array[1882]=30'd959928886;
array[1883]=30'd959928886;
array[1884]=30'd959928886;
array[1885]=30'd959928886;
array[1886]=30'd959928886;
array[1887]=30'd959928886;
array[1888]=30'd959928886;
array[1889]=30'd959928886;
array[1890]=30'd959928886;
array[1891]=30'd916921900;
array[1892]=30'd555187752;
array[1893]=30'd401043987;
array[1894]=30'd959928886;
array[1895]=30'd938933826;
array[1896]=30'd712431145;
array[1897]=30'd625322602;
array[1898]=30'd608527024;
array[1899]=30'd393597595;
array[1900]=30'd559255224;
array[1901]=30'd646262454;
array[1902]=30'd516257448;
array[1903]=30'd608527024;
array[1904]=30'd608527024;
array[1905]=30'd709306968;
array[1906]=30'd884420162;
array[1907]=30'd879168118;
array[1908]=30'd879168118;
array[1909]=30'd879168118;
array[1910]=30'd898043496;
array[1911]=30'd898043496;
array[1912]=30'd898043496;
array[1913]=30'd898043496;
array[1914]=30'd879168118;
array[1915]=30'd879168118;
array[1916]=30'd879168118;
array[1917]=30'd879168118;
array[1918]=30'd856066696;
array[1919]=30'd856066696;
array[1920]=30'd879168118;
array[1921]=30'd856066696;
array[1922]=30'd879168118;
array[1923]=30'd879168118;
array[1924]=30'd879168118;
array[1925]=30'd879168118;
array[1926]=30'd879168118;
array[1927]=30'd879168118;
array[1928]=30'd879168118;
array[1929]=30'd879168118;
array[1930]=30'd898043496;
array[1931]=30'd959928886;
array[1932]=30'd821544417;
array[1933]=30'd425179585;
array[1934]=30'd472369584;
array[1935]=30'd472369584;
array[1936]=30'd472369584;
array[1937]=30'd396870070;
array[1938]=30'd472369584;
array[1939]=30'd472369584;
array[1940]=30'd472369584;
array[1941]=30'd740803022;
array[1942]=30'd821544417;
array[1943]=30'd860309028;
array[1944]=30'd879168118;
array[1945]=30'd879168118;
array[1946]=30'd879168118;
array[1947]=30'd879168118;
array[1948]=30'd879168118;
array[1949]=30'd879168118;
array[1950]=30'd879168118;
array[1951]=30'd879168118;
array[1952]=30'd879168118;
array[1953]=30'd879168118;
array[1954]=30'd879168118;
array[1955]=30'd856066696;
array[1956]=30'd856066696;
array[1957]=30'd856066696;
array[1958]=30'd856066696;
array[1959]=30'd879168118;
array[1960]=30'd729186945;
array[1961]=30'd559255224;
array[1962]=30'd646262454;
array[1963]=30'd485848753;
array[1964]=30'd669371047;
array[1965]=30'd558250630;
array[1966]=30'd938933826;
array[1967]=30'd938933826;
array[1968]=30'd959928886;
array[1969]=30'd959928886;
array[1970]=30'd959928886;
array[1971]=30'd959928886;
array[1972]=30'd959928886;
array[1973]=30'd959928886;
array[1974]=30'd959928886;
array[1975]=30'd979842606;
array[1976]=30'd979842606;
array[1977]=30'd979842606;
array[1978]=30'd979842606;
array[1979]=30'd959928886;
array[1980]=30'd959928886;
array[1981]=30'd959928886;
array[1982]=30'd959928886;
array[1983]=30'd959928886;
array[1984]=30'd959928886;
array[1985]=30'd959928886;
array[1986]=30'd959928886;
array[1987]=30'd959928886;
array[1988]=30'd938933826;
array[1989]=30'd810005031;
array[1990]=30'd959928886;
array[1991]=30'd938933826;
array[1992]=30'd624350812;
array[1993]=30'd665151100;
array[1994]=30'd613805729;
array[1995]=30'd362130088;
array[1996]=30'd608527024;
array[1997]=30'd646262454;
array[1998]=30'd485848753;
array[1999]=30'd646262454;
array[2000]=30'd551919254;
array[2001]=30'd815194717;
array[2002]=30'd959928886;
array[2003]=30'd884420162;
array[2004]=30'd916921900;
array[2005]=30'd916921900;
array[2006]=30'd903304711;
array[2007]=30'd945268200;
array[2008]=30'd945268200;
array[2009]=30'd960978443;
array[2010]=30'd959928886;
array[2011]=30'd938933826;
array[2012]=30'd879168118;
array[2013]=30'd856066696;
array[2014]=30'd856066696;
array[2015]=30'd856066696;
array[2016]=30'd879168118;
array[2017]=30'd856066696;
array[2018]=30'd879168118;
array[2019]=30'd879168118;
array[2020]=30'd879168118;
array[2021]=30'd879168118;
array[2022]=30'd879168118;
array[2023]=30'd879168118;
array[2024]=30'd879168118;
array[2025]=30'd879168118;
array[2026]=30'd938933826;
array[2027]=30'd936883742;
array[2028]=30'd775423471;
array[2029]=30'd674763200;
array[2030]=30'd472369584;
array[2031]=30'd472369584;
array[2032]=30'd472369584;
array[2033]=30'd425179585;
array[2034]=30'd425179585;
array[2035]=30'd472369584;
array[2036]=30'd674763200;
array[2037]=30'd798493124;
array[2038]=30'd798493124;
array[2039]=30'd860309028;
array[2040]=30'd879168118;
array[2041]=30'd879168118;
array[2042]=30'd879168118;
array[2043]=30'd879168118;
array[2044]=30'd879168118;
array[2045]=30'd879168118;
array[2046]=30'd879168118;
array[2047]=30'd879168118;
array[2048]=30'd879168118;
array[2049]=30'd879168118;
array[2050]=30'd879168118;
array[2051]=30'd856066696;
array[2052]=30'd879168118;
array[2053]=30'd856066696;
array[2054]=30'd856066696;
array[2055]=30'd879168118;
array[2056]=30'd781608573;
array[2057]=30'd551919254;
array[2058]=30'd646262454;
array[2059]=30'd444952244;
array[2060]=30'd669371047;
array[2061]=30'd558250630;
array[2062]=30'd842499661;
array[2063]=30'd916921900;
array[2064]=30'd884420162;
array[2065]=30'd916921900;
array[2066]=30'd938933826;
array[2067]=30'd916921900;
array[2068]=30'd959928886;
array[2069]=30'd959928886;
array[2070]=30'd959928886;
array[2071]=30'd959928886;
array[2072]=30'd959928886;
array[2073]=30'd959928886;
array[2074]=30'd979842606;
array[2075]=30'd959928886;
array[2076]=30'd959928886;
array[2077]=30'd959928886;
array[2078]=30'd959928886;
array[2079]=30'd959928886;
array[2080]=30'd959928886;
array[2081]=30'd884420162;
array[2082]=30'd959928886;
array[2083]=30'd938933826;
array[2084]=30'd884420162;
array[2085]=30'd959928886;
array[2086]=30'd938933826;
array[2087]=30'd916921900;
array[2088]=30'd527847013;
array[2089]=30'd665151100;
array[2090]=30'd559255224;
array[2091]=30'd427157133;
array[2092]=30'd646262454;
array[2093]=30'd646262454;
array[2094]=30'd516257448;
array[2095]=30'd646262454;
array[2096]=30'd522581659;
array[2097]=30'd795279924;
array[2098]=30'd903304711;
array[2099]=30'd843548160;
array[2100]=30'd785935846;
array[2101]=30'd758671804;
array[2102]=30'd758671804;
array[2103]=30'd774396326;
array[2104]=30'd774396326;
array[2105]=30'd816348600;
array[2106]=30'd898119130;
array[2107]=30'd960978443;
array[2108]=30'd884420162;
array[2109]=30'd879168118;
array[2110]=30'd856066696;
array[2111]=30'd856066696;
array[2112]=30'd879168118;
array[2113]=30'd879168118;
array[2114]=30'd879168118;
array[2115]=30'd879168118;
array[2116]=30'd879168118;
array[2117]=30'd879168118;
array[2118]=30'd879168118;
array[2119]=30'd879168118;
array[2120]=30'd879168118;
array[2121]=30'd879168118;
array[2122]=30'd919054939;
array[2123]=30'd827871766;
array[2124]=30'd821544417;
array[2125]=30'd881300969;
array[2126]=30'd746067471;
array[2127]=30'd456626661;
array[2128]=30'd472369584;
array[2129]=30'd472369584;
array[2130]=30'd425179585;
array[2131]=30'd425179585;
array[2132]=30'd821544417;
array[2133]=30'd821544417;
array[2134]=30'd798493124;
array[2135]=30'd903304711;
array[2136]=30'd879168118;
array[2137]=30'd879168118;
array[2138]=30'd879168118;
array[2139]=30'd879168118;
array[2140]=30'd879168118;
array[2141]=30'd879168118;
array[2142]=30'd879168118;
array[2143]=30'd879168118;
array[2144]=30'd879168118;
array[2145]=30'd879168118;
array[2146]=30'd879168118;
array[2147]=30'd856066696;
array[2148]=30'd879168118;
array[2149]=30'd856066696;
array[2150]=30'd856066696;
array[2151]=30'd879168118;
array[2152]=30'd814111379;
array[2153]=30'd522581659;
array[2154]=30'd646262454;
array[2155]=30'd452327079;
array[2156]=30'd646262454;
array[2157]=30'd624350812;
array[2158]=30'd938933826;
array[2159]=30'd938933826;
array[2160]=30'd884420162;
array[2161]=30'd959928886;
array[2162]=30'd959928886;
array[2163]=30'd959928886;
array[2164]=30'd959928886;
array[2165]=30'd959928886;
array[2166]=30'd959928886;
array[2167]=30'd959928886;
array[2168]=30'd959928886;
array[2169]=30'd959928886;
array[2170]=30'd959928886;
array[2171]=30'd979842606;
array[2172]=30'd979842606;
array[2173]=30'd979842606;
array[2174]=30'd959928886;
array[2175]=30'd959928886;
array[2176]=30'd916921900;
array[2177]=30'd938933826;
array[2178]=30'd959928886;
array[2179]=30'd884420162;
array[2180]=30'd959928886;
array[2181]=30'd959928886;
array[2182]=30'd841408084;
array[2183]=30'd860309028;
array[2184]=30'd527847013;
array[2185]=30'd634745492;
array[2186]=30'd522581659;
array[2187]=30'd496374434;
array[2188]=30'd646262454;
array[2189]=30'd581260986;
array[2190]=30'd559255224;
array[2191]=30'd646262454;
array[2192]=30'd558250630;
array[2193]=30'd860309028;
array[2194]=30'd775423471;
array[2195]=30'd775423471;
array[2196]=30'd785935846;
array[2197]=30'd816348600;
array[2198]=30'd850952611;
array[2199]=30'd885566856;
array[2200]=30'd885566856;
array[2201]=30'd832088453;
array[2202]=30'd790145435;
array[2203]=30'd945268200;
array[2204]=30'd916921900;
array[2205]=30'd841408084;
array[2206]=30'd856066696;
array[2207]=30'd856066696;
array[2208]=30'd879168118;
array[2209]=30'd879168118;
array[2210]=30'd879168118;
array[2211]=30'd879168118;
array[2212]=30'd879168118;
array[2213]=30'd879168118;
array[2214]=30'd879168118;
array[2215]=30'd879168118;
array[2216]=30'd879168118;
array[2217]=30'd879168118;
array[2218]=30'd898043496;
array[2219]=30'd898098744;
array[2220]=30'd884420162;
array[2221]=30'd884420162;
array[2222]=30'd884420162;
array[2223]=30'd725052963;
array[2224]=30'd463997419;
array[2225]=30'd472369584;
array[2226]=30'd472369584;
array[2227]=30'd425179585;
array[2228]=30'd843548160;
array[2229]=30'd903304711;
array[2230]=30'd903304711;
array[2231]=30'd860309028;
array[2232]=30'd879168118;
array[2233]=30'd879168118;
array[2234]=30'd879168118;
array[2235]=30'd879168118;
array[2236]=30'd879168118;
array[2237]=30'd879168118;
array[2238]=30'd879168118;
array[2239]=30'd879168118;
array[2240]=30'd879168118;
array[2241]=30'd879168118;
array[2242]=30'd879168118;
array[2243]=30'd879168118;
array[2244]=30'd879168118;
array[2245]=30'd879168118;
array[2246]=30'd879168118;
array[2247]=30'd879168118;
array[2248]=30'd856066696;
array[2249]=30'd558250630;
array[2250]=30'd634745492;
array[2251]=30'd452327079;
array[2252]=30'd613805729;
array[2253]=30'd729186945;
array[2254]=30'd959928886;
array[2255]=30'd959928886;
array[2256]=30'd959928886;
array[2257]=30'd959928886;
array[2258]=30'd959928886;
array[2259]=30'd959928886;
array[2260]=30'd959928886;
array[2261]=30'd959928886;
array[2262]=30'd959928886;
array[2263]=30'd959928886;
array[2264]=30'd959928886;
array[2265]=30'd959928886;
array[2266]=30'd959928886;
array[2267]=30'd959928886;
array[2268]=30'd959928886;
array[2269]=30'd959928886;
array[2270]=30'd959928886;
array[2271]=30'd959928886;
array[2272]=30'd959928886;
array[2273]=30'd959928886;
array[2274]=30'd959928886;
array[2275]=30'd959928886;
array[2276]=30'd959928886;
array[2277]=30'd938933826;
array[2278]=30'd938933826;
array[2279]=30'd795279924;
array[2280]=30'd582343294;
array[2281]=30'd634745492;
array[2282]=30'd467006094;
array[2283]=30'd559255224;
array[2284]=30'd646262454;
array[2285]=30'd516257448;
array[2286]=30'd581260986;
array[2287]=30'd608527024;
array[2288]=30'd641178190;
array[2289]=30'd827871766;
array[2290]=30'd798493124;
array[2291]=30'd871910847;
array[2292]=30'd898119130;
array[2293]=30'd871910847;
array[2294]=30'd871910847;
array[2295]=30'd850952611;
array[2296]=30'd850952611;
array[2297]=30'd850952611;
array[2298]=30'd790145435;
array[2299]=30'd871910847;
array[2300]=30'd960978443;
array[2301]=30'd884420162;
array[2302]=30'd879168118;
array[2303]=30'd856066696;
array[2304]=30'd898043496;
array[2305]=30'd898043496;
array[2306]=30'd879168118;
array[2307]=30'd879168118;
array[2308]=30'd879168118;
array[2309]=30'd879168118;
array[2310]=30'd879168118;
array[2311]=30'd898043496;
array[2312]=30'd879168118;
array[2313]=30'd879168118;
array[2314]=30'd879168118;
array[2315]=30'd898043496;
array[2316]=30'd879168118;
array[2317]=30'd898043496;
array[2318]=30'd879168118;
array[2319]=30'd898043496;
array[2320]=30'd725052963;
array[2321]=30'd456626661;
array[2322]=30'd472369584;
array[2323]=30'd425179585;
array[2324]=30'd725052963;
array[2325]=30'd884420162;
array[2326]=30'd884420162;
array[2327]=30'd879168118;
array[2328]=30'd879168118;
array[2329]=30'd879168118;
array[2330]=30'd879168118;
array[2331]=30'd879168118;
array[2332]=30'd879168118;
array[2333]=30'd879168118;
array[2334]=30'd879168118;
array[2335]=30'd879168118;
array[2336]=30'd879168118;
array[2337]=30'd879168118;
array[2338]=30'd879168118;
array[2339]=30'd879168118;
array[2340]=30'd879168118;
array[2341]=30'd879168118;
array[2342]=30'd879168118;
array[2343]=30'd879168118;
array[2344]=30'd856066696;
array[2345]=30'd605405812;
array[2346]=30'd634745492;
array[2347]=30'd467006094;
array[2348]=30'd559255224;
array[2349]=30'd815194717;
array[2350]=30'd979842606;
array[2351]=30'd959928886;
array[2352]=30'd959928886;
array[2353]=30'd959928886;
array[2354]=30'd959928886;
array[2355]=30'd668430907;
array[2356]=30'd597116464;
array[2357]=30'd641178190;
array[2358]=30'd694642226;
array[2359]=30'd756500033;
array[2360]=30'd795279924;
array[2361]=30'd810005031;
array[2362]=30'd795279924;
array[2363]=30'd795279924;
array[2364]=30'd756500033;
array[2365]=30'd725052963;
array[2366]=30'd668430907;
array[2367]=30'd612873765;
array[2368]=30'd528973367;
array[2369]=30'd668430907;
array[2370]=30'd959928886;
array[2371]=30'd959928886;
array[2372]=30'd959928886;
array[2373]=30'd959928886;
array[2374]=30'd938933826;
array[2375]=30'd709306968;
array[2376]=30'd605405812;
array[2377]=30'd608527024;
array[2378]=30'd427157133;
array[2379]=30'd608527024;
array[2380]=30'd608527024;
array[2381]=30'd467006094;
array[2382]=30'd608527024;
array[2383]=30'd551919254;
array[2384]=30'd709306968;
array[2385]=30'd785935846;
array[2386]=30'd833115609;
array[2387]=30'd925360587;
array[2388]=30'd833115609;
array[2389]=30'd758671804;
array[2390]=30'd758671804;
array[2391]=30'd774396326;
array[2392]=30'd763929993;
array[2393]=30'd790145435;
array[2394]=30'd832088453;
array[2395]=30'd816348600;
array[2396]=30'd945268200;
array[2397]=30'd916921900;
array[2398]=30'd879168118;
array[2399]=30'd856066696;
array[2400]=30'd884420162;
array[2401]=30'd860309028;
array[2402]=30'd884420162;
array[2403]=30'd884420162;
array[2404]=30'd898043496;
array[2405]=30'd898043496;
array[2406]=30'd879168118;
array[2407]=30'd879168118;
array[2408]=30'd879168118;
array[2409]=30'd898043496;
array[2410]=30'd898043496;
array[2411]=30'd898043496;
array[2412]=30'd879168118;
array[2413]=30'd879168118;
array[2414]=30'd879168118;
array[2415]=30'd879168118;
array[2416]=30'd884420162;
array[2417]=30'd475488805;
array[2418]=30'd484957641;
array[2419]=30'd477594065;
array[2420]=30'd617030138;
array[2421]=30'd884420162;
array[2422]=30'd879168118;
array[2423]=30'd879168118;
array[2424]=30'd879168118;
array[2425]=30'd879168118;
array[2426]=30'd879168118;
array[2427]=30'd879168118;
array[2428]=30'd879168118;
array[2429]=30'd879168118;
array[2430]=30'd879168118;
array[2431]=30'd879168118;
array[2432]=30'd879168118;
array[2433]=30'd879168118;
array[2434]=30'd879168118;
array[2435]=30'd879168118;
array[2436]=30'd879168118;
array[2437]=30'd879168118;
array[2438]=30'd879168118;
array[2439]=30'd879168118;
array[2440]=30'd879168118;
array[2441]=30'd686214797;
array[2442]=30'd582343294;
array[2443]=30'd427157133;
array[2444]=30'd582343294;
array[2445]=30'd815194717;
array[2446]=30'd959928886;
array[2447]=30'd959928886;
array[2448]=30'd959928886;
array[2449]=30'd959928886;
array[2450]=30'd959928886;
array[2451]=30'd612873765;
array[2452]=30'd377963103;
array[2453]=30'd377963103;
array[2454]=30'd377963103;
array[2455]=30'd377963103;
array[2456]=30'd377963103;
array[2457]=30'd377963103;
array[2458]=30'd377963103;
array[2459]=30'd377963103;
array[2460]=30'd377963103;
array[2461]=30'd377963103;
array[2462]=30'd377963103;
array[2463]=30'd377963103;
array[2464]=30'd377963103;
array[2465]=30'd475488805;
array[2466]=30'd959928886;
array[2467]=30'd959928886;
array[2468]=30'd959928886;
array[2469]=30'd959928886;
array[2470]=30'd938933826;
array[2471]=30'd624350812;
array[2472]=30'd634745492;
array[2473]=30'd613805729;
array[2474]=30'd496374434;
array[2475]=30'd634745492;
array[2476]=30'd559255224;
array[2477]=30'd427157133;
array[2478]=30'd634745492;
array[2479]=30'd558250630;
array[2480]=30'd779606588;
array[2481]=30'd758671804;
array[2482]=30'd871910847;
array[2483]=30'd881300969;
array[2484]=30'd785935846;
array[2485]=30'd758671804;
array[2486]=30'd911766951;
array[2487]=30'd871910847;
array[2488]=30'd790145435;
array[2489]=30'd790145435;
array[2490]=30'd885566856;
array[2491]=30'd790145435;
array[2492]=30'd925360587;
array[2493]=30'd936883742;
array[2494]=30'd884420162;
array[2495]=30'd879168118;
array[2496]=30'd843548160;
array[2497]=30'd843548160;
array[2498]=30'd843548160;
array[2499]=30'd903304711;
array[2500]=30'd884420162;
array[2501]=30'd898043496;
array[2502]=30'd879168118;
array[2503]=30'd879168118;
array[2504]=30'd879168118;
array[2505]=30'd879168118;
array[2506]=30'd898043496;
array[2507]=30'd898043496;
array[2508]=30'd898043496;
array[2509]=30'd898043496;
array[2510]=30'd898043496;
array[2511]=30'd879168118;
array[2512]=30'd879168118;
array[2513]=30'd597116464;
array[2514]=30'd484957641;
array[2515]=30'd477594065;
array[2516]=30'd515315216;
array[2517]=30'd884420162;
array[2518]=30'd879168118;
array[2519]=30'd879168118;
array[2520]=30'd898043496;
array[2521]=30'd879168118;
array[2522]=30'd879168118;
array[2523]=30'd898043496;
array[2524]=30'd879168118;
array[2525]=30'd879168118;
array[2526]=30'd879168118;
array[2527]=30'd879168118;
array[2528]=30'd879168118;
array[2529]=30'd879168118;
array[2530]=30'd879168118;
array[2531]=30'd879168118;
array[2532]=30'd879168118;
array[2533]=30'd879168118;
array[2534]=30'd879168118;
array[2535]=30'd879168118;
array[2536]=30'd879168118;
array[2537]=30'd781608573;
array[2538]=30'd527847013;
array[2539]=30'd427157133;
array[2540]=30'd669371047;
array[2541]=30'd683036269;
array[2542]=30'd959928886;
array[2543]=30'd959928886;
array[2544]=30'd959928886;
array[2545]=30'd959928886;
array[2546]=30'd959928886;
array[2547]=30'd756500033;
array[2548]=30'd344392301;
array[2549]=30'd398924382;
array[2550]=30'd398924382;
array[2551]=30'd398924382;
array[2552]=30'd398924382;
array[2553]=30'd398924382;
array[2554]=30'd398924382;
array[2555]=30'd377963103;
array[2556]=30'd377963103;
array[2557]=30'd377963103;
array[2558]=30'd398924382;
array[2559]=30'd398924382;
array[2560]=30'd377963103;
array[2561]=30'd571952708;
array[2562]=30'd959928886;
array[2563]=30'd959928886;
array[2564]=30'd959928886;
array[2565]=30'd938933826;
array[2566]=30'd916921900;
array[2567]=30'd559303250;
array[2568]=30'd634745492;
array[2569]=30'd551919254;
array[2570]=30'd581260986;
array[2571]=30'd608527024;
array[2572]=30'd427157133;
array[2573]=30'd522581659;
array[2574]=30'd634745492;
array[2575]=30'd566698607;
array[2576]=30'd810005031;
array[2577]=30'd816348600;
array[2578]=30'd925360587;
array[2579]=30'd881300969;
array[2580]=30'd785935846;
array[2581]=30'd816348600;
array[2582]=30'd945316283;
array[2583]=30'd911766951;
array[2584]=30'd816348600;
array[2585]=30'd790145435;
array[2586]=30'd911766951;
array[2587]=30'd790145435;
array[2588]=30'd871910847;
array[2589]=30'd903304711;
array[2590]=30'd884420162;
array[2591]=30'd879168118;
array[2592]=30'd857224695;
array[2593]=30'd852996553;
array[2594]=30'd881300969;
array[2595]=30'd903304711;
array[2596]=30'd884420162;
array[2597]=30'd898043496;
array[2598]=30'd879168118;
array[2599]=30'd898043496;
array[2600]=30'd898043496;
array[2601]=30'd898043496;
array[2602]=30'd898043496;
array[2603]=30'd898043496;
array[2604]=30'd898043496;
array[2605]=30'd898043496;
array[2606]=30'd898043496;
array[2607]=30'd898043496;
array[2608]=30'd898043496;
array[2609]=30'd694642226;
array[2610]=30'd463997419;
array[2611]=30'd484957641;
array[2612]=30'd456626661;
array[2613]=30'd860309028;
array[2614]=30'd898043496;
array[2615]=30'd898043496;
array[2616]=30'd879168118;
array[2617]=30'd879168118;
array[2618]=30'd898043496;
array[2619]=30'd898043496;
array[2620]=30'd898043496;
array[2621]=30'd879168118;
array[2622]=30'd879168118;
array[2623]=30'd879168118;
array[2624]=30'd879168118;
array[2625]=30'd879168118;
array[2626]=30'd879168118;
array[2627]=30'd879168118;
array[2628]=30'd879168118;
array[2629]=30'd879168118;
array[2630]=30'd879168118;
array[2631]=30'd879168118;
array[2632]=30'd879168118;
array[2633]=30'd856066696;
array[2634]=30'd527847013;
array[2635]=30'd485876339;
array[2636]=30'd669371047;
array[2637]=30'd613805729;
array[2638]=30'd815194717;
array[2639]=30'd959928886;
array[2640]=30'd959928886;
array[2641]=30'd959928886;
array[2642]=30'd959928886;
array[2643]=30'd916921900;
array[2644]=30'd475488805;
array[2645]=30'd398924382;
array[2646]=30'd398924382;
array[2647]=30'd459725411;
array[2648]=30'd459725411;
array[2649]=30'd459725411;
array[2650]=30'd459725411;
array[2651]=30'd459725411;
array[2652]=30'd398924382;
array[2653]=30'd398924382;
array[2654]=30'd398924382;
array[2655]=30'd398924382;
array[2656]=30'd428280389;
array[2657]=30'd860309028;
array[2658]=30'd959928886;
array[2659]=30'd959928886;
array[2660]=30'd959928886;
array[2661]=30'd938933826;
array[2662]=30'd841408084;
array[2663]=30'd527847013;
array[2664]=30'd634745492;
array[2665]=30'd496374434;
array[2666]=30'd646262454;
array[2667]=30'd559255224;
array[2668]=30'd331722417;
array[2669]=30'd559255224;
array[2670]=30'd634745492;
array[2671]=30'd592910950;
array[2672]=30'd775423471;
array[2673]=30'd833115609;
array[2674]=30'd945268200;
array[2675]=30'd860309028;
array[2676]=30'd827871766;
array[2677]=30'd774396326;
array[2678]=30'd911766951;
array[2679]=30'd816348600;
array[2680]=30'd774396326;
array[2681]=30'd790145435;
array[2682]=30'd885566856;
array[2683]=30'd790145435;
array[2684]=30'd852996553;
array[2685]=30'd903304711;
array[2686]=30'd884420162;
array[2687]=30'd879168118;
array[2688]=30'd857224695;
array[2689]=30'd881300969;
array[2690]=30'd881300969;
array[2691]=30'd860309028;
array[2692]=30'd884420162;
array[2693]=30'd898043496;
array[2694]=30'd898043496;
array[2695]=30'd898043496;
array[2696]=30'd898043496;
array[2697]=30'd898043496;
array[2698]=30'd898043496;
array[2699]=30'd898043496;
array[2700]=30'd898043496;
array[2701]=30'd898043496;
array[2702]=30'd898043496;
array[2703]=30'd898043496;
array[2704]=30'd898043496;
array[2705]=30'd799523423;
array[2706]=30'd596111858;
array[2707]=30'd775423471;
array[2708]=30'd843548160;
array[2709]=30'd756500033;
array[2710]=30'd898043496;
array[2711]=30'd898043496;
array[2712]=30'd898043496;
array[2713]=30'd898043496;
array[2714]=30'd898043496;
array[2715]=30'd898043496;
array[2716]=30'd898043496;
array[2717]=30'd898043496;
array[2718]=30'd898043496;
array[2719]=30'd898043496;
array[2720]=30'd898043496;
array[2721]=30'd898043496;
array[2722]=30'd898043496;
array[2723]=30'd879168118;
array[2724]=30'd879168118;
array[2725]=30'd879168118;
array[2726]=30'd879168118;
array[2727]=30'd879168118;
array[2728]=30'd879168118;
array[2729]=30'd879168118;
array[2730]=30'd527847013;
array[2731]=30'd448143984;
array[2732]=30'd646262454;
array[2733]=30'd608527024;
array[2734]=30'd483822211;
array[2735]=30'd709306968;
array[2736]=30'd959928886;
array[2737]=30'd959928886;
array[2738]=30'd959928886;
array[2739]=30'd959928886;
array[2740]=30'd884420162;
array[2741]=30'd548890196;
array[2742]=30'd571952708;
array[2743]=30'd624350812;
array[2744]=30'd624350812;
array[2745]=30'd624350812;
array[2746]=30'd624350812;
array[2747]=30'd624350812;
array[2748]=30'd592910950;
array[2749]=30'd530016882;
array[2750]=30'd459725411;
array[2751]=30'd428280389;
array[2752]=30'd795279924;
array[2753]=30'd959928886;
array[2754]=30'd959928886;
array[2755]=30'd959928886;
array[2756]=30'd938933826;
array[2757]=30'd938933826;
array[2758]=30'd665233987;
array[2759]=30'd582343294;
array[2760]=30'd551919254;
array[2761]=30'd559255224;
array[2762]=30'd608527024;
array[2763]=30'd452327079;
array[2764]=30'd393597595;
array[2765]=30'd613805729;
array[2766]=30'd605405812;
array[2767]=30'd641178190;
array[2768]=30'd775423471;
array[2769]=30'd833115609;
array[2770]=30'd945268200;
array[2771]=30'd877139478;
array[2772]=30'd785935846;
array[2773]=30'd758671804;
array[2774]=30'd945316283;
array[2775]=30'd871910847;
array[2776]=30'd816348600;
array[2777]=30'd816348600;
array[2778]=30'd790145435;
array[2779]=30'd774396326;
array[2780]=30'd881300969;
array[2781]=30'd860309028;
array[2782]=30'd879168118;
array[2783]=30'd879168118;
array[2784]=30'd877139478;
array[2785]=30'd877139478;
array[2786]=30'd903304711;
array[2787]=30'd884420162;
array[2788]=30'd898043496;
array[2789]=30'd898043496;
array[2790]=30'd898043496;
array[2791]=30'd898043496;
array[2792]=30'd898043496;
array[2793]=30'd879168118;
array[2794]=30'd898043496;
array[2795]=30'd898043496;
array[2796]=30'd898043496;
array[2797]=30'd898043496;
array[2798]=30'd898043496;
array[2799]=30'd898043496;
array[2800]=30'd898043496;
array[2801]=30'd884420162;
array[2802]=30'd810005031;
array[2803]=30'd1034407430;
array[2804]=30'd960978443;
array[2805]=30'd712431145;
array[2806]=30'd898043496;
array[2807]=30'd898043496;
array[2808]=30'd898043496;
array[2809]=30'd898043496;
array[2810]=30'd898043496;
array[2811]=30'd898043496;
array[2812]=30'd898043496;
array[2813]=30'd898043496;
array[2814]=30'd898043496;
array[2815]=30'd898043496;
array[2816]=30'd898043496;
array[2817]=30'd898043496;
array[2818]=30'd898043496;
array[2819]=30'd898043496;
array[2820]=30'd898043496;
array[2821]=30'd898043496;
array[2822]=30'd898043496;
array[2823]=30'd898043496;
array[2824]=30'd879168118;
array[2825]=30'd879168118;
array[2826]=30'd624350812;
array[2827]=30'd448143984;
array[2828]=30'd646262454;
array[2829]=30'd608527024;
array[2830]=30'd452327079;
array[2831]=30'd434534016;
array[2832]=30'd624350812;
array[2833]=30'd884420162;
array[2834]=30'd959928886;
array[2835]=30'd959928886;
array[2836]=30'd938933826;
array[2837]=30'd916921900;
array[2838]=30'd756500033;
array[2839]=30'd571952708;
array[2840]=30'd548890196;
array[2841]=30'd548890196;
array[2842]=30'd566698607;
array[2843]=30'd548890196;
array[2844]=30'd548890196;
array[2845]=30'd548890196;
array[2846]=30'd709306968;
array[2847]=30'd884420162;
array[2848]=30'd959928886;
array[2849]=30'd959928886;
array[2850]=30'd959928886;
array[2851]=30'd959928886;
array[2852]=30'd884420162;
array[2853]=30'd597116464;
array[2854]=30'd361121389;
array[2855]=30'd634745492;
array[2856]=30'd452327079;
array[2857]=30'd608527024;
array[2858]=30'd551919254;
array[2859]=30'd331722417;
array[2860]=30'd467006094;
array[2861]=30'd634745492;
array[2862]=30'd582343294;
array[2863]=30'd744990312;
array[2864]=30'd746067471;
array[2865]=30'd833115609;
array[2866]=30'd964180446;
array[2867]=30'd936883742;
array[2868]=30'd827871766;
array[2869]=30'd758671804;
array[2870]=30'd911766951;
array[2871]=30'd977825191;
array[2872]=30'd945316283;
array[2873]=30'd911766951;
array[2874]=30'd774396326;
array[2875]=30'd852996553;
array[2876]=30'd903304711;
array[2877]=30'd884420162;
array[2878]=30'd879168118;
array[2879]=30'd879168118;
array[2880]=30'd877139478;
array[2881]=30'd877139478;
array[2882]=30'd884420162;
array[2883]=30'd884420162;
array[2884]=30'd898043496;
array[2885]=30'd898043496;
array[2886]=30'd898043496;
array[2887]=30'd898043496;
array[2888]=30'd898043496;
array[2889]=30'd898043496;
array[2890]=30'd898043496;
array[2891]=30'd898043496;
array[2892]=30'd879168118;
array[2893]=30'd898043496;
array[2894]=30'd879168118;
array[2895]=30'd879168118;
array[2896]=30'd898043496;
array[2897]=30'd898043496;
array[2898]=30'd756500033;
array[2899]=30'd1034407430;
array[2900]=30'd1000848926;
array[2901]=30'd725052963;
array[2902]=30'd898043496;
array[2903]=30'd898043496;
array[2904]=30'd898043496;
array[2905]=30'd898043496;
array[2906]=30'd898043496;
array[2907]=30'd898043496;
array[2908]=30'd898043496;
array[2909]=30'd898043496;
array[2910]=30'd898043496;
array[2911]=30'd898043496;
array[2912]=30'd884420162;
array[2913]=30'd884420162;
array[2914]=30'd898043496;
array[2915]=30'd898043496;
array[2916]=30'd898043496;
array[2917]=30'd898043496;
array[2918]=30'd898043496;
array[2919]=30'd898043496;
array[2920]=30'd879168118;
array[2921]=30'd879168118;
array[2922]=30'd709306968;
array[2923]=30'd485876339;
array[2924]=30'd634745492;
array[2925]=30'd559255224;
array[2926]=30'd452327079;
array[2927]=30'd467006094;
array[2928]=30'd361121389;
array[2929]=30'd459725411;
array[2930]=30'd709306968;
array[2931]=30'd916921900;
array[2932]=30'd959928886;
array[2933]=30'd959928886;
array[2934]=30'd959928886;
array[2935]=30'd959928886;
array[2936]=30'd884420162;
array[2937]=30'd860309028;
array[2938]=30'd860309028;
array[2939]=30'd884420162;
array[2940]=30'd916921900;
array[2941]=30'd959928886;
array[2942]=30'd959928886;
array[2943]=30'd959928886;
array[2944]=30'd959928886;
array[2945]=30'd959928886;
array[2946]=30'd938933826;
array[2947]=30'd756500033;
array[2948]=30'd462859830;
array[2949]=30'd414594647;
array[2950]=30'd448143984;
array[2951]=30'd582343294;
array[2952]=30'd516257448;
array[2953]=30'd608527024;
array[2954]=30'd393597595;
array[2955]=30'd340142721;
array[2956]=30'd467006094;
array[2957]=30'd634745492;
array[2958]=30'd551919254;
array[2959]=30'd799523423;
array[2960]=30'd827871766;
array[2961]=30'd798493124;
array[2962]=30'd945316283;
array[2963]=30'd983039487;
array[2964]=30'd877139478;
array[2965]=30'd785935846;
array[2966]=30'd774396326;
array[2967]=30'd850952611;
array[2968]=30'd871910847;
array[2969]=30'd816348600;
array[2970]=30'd774396326;
array[2971]=30'd881300969;
array[2972]=30'd903304711;
array[2973]=30'd898043496;
array[2974]=30'd898043496;
array[2975]=30'd879168118;
array[2976]=30'd884420162;
array[2977]=30'd884420162;
array[2978]=30'd884420162;
array[2979]=30'd898043496;
array[2980]=30'd898043496;
array[2981]=30'd879168118;
array[2982]=30'd898043496;
array[2983]=30'd898043496;
array[2984]=30'd898043496;
array[2985]=30'd898043496;
array[2986]=30'd898043496;
array[2987]=30'd898043496;
array[2988]=30'd879168118;
array[2989]=30'd898043496;
array[2990]=30'd898043496;
array[2991]=30'd898043496;
array[2992]=30'd898043496;
array[2993]=30'd898043496;
array[2994]=30'd725091917;
array[2995]=30'd1034407430;
array[2996]=30'd1034407430;
array[2997]=30'd795279924;
array[2998]=30'd884420162;
array[2999]=30'd898043496;
array[3000]=30'd898043496;
array[3001]=30'd898043496;
array[3002]=30'd898043496;
array[3003]=30'd898043496;
array[3004]=30'd898043496;
array[3005]=30'd898043496;
array[3006]=30'd898043496;
array[3007]=30'd898043496;
array[3008]=30'd810005031;
array[3009]=30'd936883742;
array[3010]=30'd898098744;
array[3011]=30'd860309028;
array[3012]=30'd916921900;
array[3013]=30'd898043496;
array[3014]=30'd898043496;
array[3015]=30'd879168118;
array[3016]=30'd879168118;
array[3017]=30'd879168118;
array[3018]=30'd739680847;
array[3019]=30'd527847013;
array[3020]=30'd634745492;
array[3021]=30'd559255224;
array[3022]=30'd452327079;
array[3023]=30'd427157133;
array[3024]=30'd340142721;
array[3025]=30'd448143984;
array[3026]=30'd414594647;
array[3027]=30'd398924382;
array[3028]=30'd624350812;
array[3029]=30'd795279924;
array[3030]=30'd916921900;
array[3031]=30'd938933826;
array[3032]=30'd959928886;
array[3033]=30'd959928886;
array[3034]=30'd959928886;
array[3035]=30'd959928886;
array[3036]=30'd959928886;
array[3037]=30'd959928886;
array[3038]=30'd959928886;
array[3039]=30'd959928886;
array[3040]=30'd884420162;
array[3041]=30'd756500033;
array[3042]=30'd512140869;
array[3043]=30'd428280389;
array[3044]=30'd448143984;
array[3045]=30'd387329638;
array[3046]=30'd527847013;
array[3047]=30'd467006094;
array[3048]=30'd613805729;
array[3049]=30'd496374434;
array[3050]=30'd281408163;
array[3051]=30'd288811658;
array[3052]=30'd483822211;
array[3053]=30'd634745492;
array[3054]=30'd558250630;
array[3055]=30'd879168118;
array[3056]=30'd855119431;
array[3057]=30'd785935846;
array[3058]=30'd816348600;
array[3059]=30'd964180446;
array[3060]=30'd983039487;
array[3061]=30'd857224695;
array[3062]=30'd833115609;
array[3063]=30'd785935846;
array[3064]=30'd758671804;
array[3065]=30'd798493124;
array[3066]=30'd852996553;
array[3067]=30'd903304711;
array[3068]=30'd884420162;
array[3069]=30'd898043496;
array[3070]=30'd879168118;
array[3071]=30'd879168118;
array[3072]=30'd898043496;
array[3073]=30'd898043496;
array[3074]=30'd898043496;
array[3075]=30'd898043496;
array[3076]=30'd898043496;
array[3077]=30'd879168118;
array[3078]=30'd898043496;
array[3079]=30'd898043496;
array[3080]=30'd898043496;
array[3081]=30'd898043496;
array[3082]=30'd898043496;
array[3083]=30'd898043496;
array[3084]=30'd898043496;
array[3085]=30'd898043496;
array[3086]=30'd898043496;
array[3087]=30'd898043496;
array[3088]=30'd898043496;
array[3089]=30'd898043496;
array[3090]=30'd725091917;
array[3091]=30'd1000848926;
array[3092]=30'd1034407430;
array[3093]=30'd903304711;
array[3094]=30'd815194717;
array[3095]=30'd898043496;
array[3096]=30'd898043496;
array[3097]=30'd898043496;
array[3098]=30'd898043496;
array[3099]=30'd898043496;
array[3100]=30'd898043496;
array[3101]=30'd898043496;
array[3102]=30'd898043496;
array[3103]=30'd919054939;
array[3104]=30'd810005031;
array[3105]=30'd960978443;
array[3106]=30'd877139478;
array[3107]=30'd810005031;
array[3108]=30'd960978443;
array[3109]=30'd916921900;
array[3110]=30'd884420162;
array[3111]=30'd898043496;
array[3112]=30'd898043496;
array[3113]=30'd879168118;
array[3114]=30'd794241637;
array[3115]=30'd558250630;
array[3116]=30'd634745492;
array[3117]=30'd516257448;
array[3118]=30'd452327079;
array[3119]=30'd434534016;
array[3120]=30'd387329638;
array[3121]=30'd448143984;
array[3122]=30'd408333955;
array[3123]=30'd387329638;
array[3124]=30'd448143984;
array[3125]=30'd414594647;
array[3126]=30'd414594647;
array[3127]=30'd548890196;
array[3128]=30'd665233987;
array[3129]=30'd795279924;
array[3130]=30'd860309028;
array[3131]=30'd884420162;
array[3132]=30'd860309028;
array[3133]=30'd795279924;
array[3134]=30'd709306968;
array[3135]=30'd665233987;
array[3136]=30'd668430907;
array[3137]=30'd756500033;
array[3138]=30'd341225034;
array[3139]=30'd428280389;
array[3140]=30'd448143984;
array[3141]=30'd387329638;
array[3142]=30'd522581659;
array[3143]=30'd522581659;
array[3144]=30'd559255224;
array[3145]=30'd408333955;
array[3146]=30'd281408163;
array[3147]=30'd340142721;
array[3148]=30'd527847013;
array[3149]=30'd634745492;
array[3150]=30'd605405812;
array[3151]=30'd898043496;
array[3152]=30'd884420162;
array[3153]=30'd827871766;
array[3154]=30'd785935846;
array[3155]=30'd898119130;
array[3156]=30'd983039487;
array[3157]=30'd936883742;
array[3158]=30'd877139478;
array[3159]=30'd877139478;
array[3160]=30'd857224695;
array[3161]=30'd903304711;
array[3162]=30'd916921900;
array[3163]=30'd898043496;
array[3164]=30'd879168118;
array[3165]=30'd879168118;
array[3166]=30'd879168118;
array[3167]=30'd879168118;
array[3168]=30'd898043496;
array[3169]=30'd898043496;
array[3170]=30'd898043496;
array[3171]=30'd898043496;
array[3172]=30'd898043496;
array[3173]=30'd898043496;
array[3174]=30'd898043496;
array[3175]=30'd884420162;
array[3176]=30'd855119431;
array[3177]=30'd860309028;
array[3178]=30'd860309028;
array[3179]=30'd884420162;
array[3180]=30'd884420162;
array[3181]=30'd898043496;
array[3182]=30'd898043496;
array[3183]=30'd898043496;
array[3184]=30'd898043496;
array[3185]=30'd898043496;
array[3186]=30'd744990312;
array[3187]=30'd936883742;
array[3188]=30'd1034407430;
array[3189]=30'd936883742;
array[3190]=30'd756500033;
array[3191]=30'd898043496;
array[3192]=30'd898043496;
array[3193]=30'd898043496;
array[3194]=30'd898043496;
array[3195]=30'd898043496;
array[3196]=30'd898043496;
array[3197]=30'd898043496;
array[3198]=30'd898043496;
array[3199]=30'd919054939;
array[3200]=30'd877139478;
array[3201]=30'd936883742;
array[3202]=30'd877139478;
array[3203]=30'd857224695;
array[3204]=30'd983039487;
array[3205]=30'd903304711;
array[3206]=30'd810005031;
array[3207]=30'd884420162;
array[3208]=30'd938933826;
array[3209]=30'd879168118;
array[3210]=30'd729186945;
array[3211]=30'd582343294;
array[3212]=30'd608527024;
array[3213]=30'd485848753;
array[3214]=30'd452327079;
array[3215]=30'd408333955;
array[3216]=30'd408333955;
array[3217]=30'd427157133;
array[3218]=30'd408333955;
array[3219]=30'd361121389;
array[3220]=30'd434534016;
array[3221]=30'd427157133;
array[3222]=30'd434534016;
array[3223]=30'd448143984;
array[3224]=30'd398924382;
array[3225]=30'd459725411;
array[3226]=30'd756500033;
array[3227]=30'd795279924;
array[3228]=30'd795279924;
array[3229]=30'd794241637;
array[3230]=30'd794241637;
array[3231]=30'd815194717;
array[3232]=30'd815194717;
array[3233]=30'd756500033;
array[3234]=30'd283619908;
array[3235]=30'd323442246;
array[3236]=30'd414594647;
array[3237]=30'd434534016;
array[3238]=30'd467006094;
array[3239]=30'd559255224;
array[3240]=30'd452327079;
array[3241]=30'd288811658;
array[3242]=30'd387329638;
array[3243]=30'd361121389;
array[3244]=30'd522581659;
array[3245]=30'd608527024;
array[3246]=30'd624350812;
array[3247]=30'd898043496;
array[3248]=30'd898043496;
array[3249]=30'd898098744;
array[3250]=30'd785935846;
array[3251]=30'd785935846;
array[3252]=30'd945316283;
array[3253]=30'd1016593896;
array[3254]=30'd983039487;
array[3255]=30'd936883742;
array[3256]=30'd945268200;
array[3257]=30'd960978443;
array[3258]=30'd916921900;
array[3259]=30'd898043496;
array[3260]=30'd879168118;
array[3261]=30'd879168118;
array[3262]=30'd879168118;
array[3263]=30'd879168118;
array[3264]=30'd898043496;
array[3265]=30'd898043496;
array[3266]=30'd898043496;
array[3267]=30'd898043496;
array[3268]=30'd898043496;
array[3269]=30'd898043496;
array[3270]=30'd884420162;
array[3271]=30'd810005031;
array[3272]=30'd821544417;
array[3273]=30'd833115609;
array[3274]=30'd833115609;
array[3275]=30'd775423471;
array[3276]=30'd843548160;
array[3277]=30'd916921900;
array[3278]=30'd898043496;
array[3279]=30'd898043496;
array[3280]=30'd898043496;
array[3281]=30'd898043496;
array[3282]=30'd799523423;
array[3283]=30'd877139478;
array[3284]=30'd1034407430;
array[3285]=30'd1000848926;
array[3286]=30'd725052963;
array[3287]=30'd938933826;
array[3288]=30'd898043496;
array[3289]=30'd898043496;
array[3290]=30'd898043496;
array[3291]=30'd898043496;
array[3292]=30'd898043496;
array[3293]=30'd898043496;
array[3294]=30'd898043496;
array[3295]=30'd919054939;
array[3296]=30'd898098744;
array[3297]=30'd898098744;
array[3298]=30'd877139478;
array[3299]=30'd921177592;
array[3300]=30'd936883742;
array[3301]=30'd843548160;
array[3302]=30'd921177592;
array[3303]=30'd960978443;
array[3304]=30'd898043496;
array[3305]=30'd879168118;
array[3306]=30'd729186945;
array[3307]=30'd634745492;
array[3308]=30'd608527024;
array[3309]=30'd444952244;
array[3310]=30'd427157133;
array[3311]=30'd344392301;
array[3312]=30'd387329638;
array[3313]=30'd448143984;
array[3314]=30'd408333955;
array[3315]=30'd289838696;
array[3316]=30'd448143984;
array[3317]=30'd448143984;
array[3318]=30'd427157133;
array[3319]=30'd434534016;
array[3320]=30'd344392301;
array[3321]=30'd344392301;
array[3322]=30'd815194717;
array[3323]=30'd815194717;
array[3324]=30'd815194717;
array[3325]=30'd815194717;
array[3326]=30'd815194717;
array[3327]=30'd815194717;
array[3328]=30'd668430907;
array[3329]=30'd428280389;
array[3330]=30'd259510865;
array[3331]=30'd283619908;
array[3332]=30'd267838034;
array[3333]=30'd448143984;
array[3334]=30'd522581659;
array[3335]=30'd516257448;
array[3336]=30'd362130088;
array[3337]=30'd344392301;
array[3338]=30'd387329638;
array[3339]=30'd361121389;
array[3340]=30'd522581659;
array[3341]=30'd613805729;
array[3342]=30'd683036269;
array[3343]=30'd898043496;
array[3344]=30'd898043496;
array[3345]=30'd919054939;
array[3346]=30'd877139478;
array[3347]=30'd785935846;
array[3348]=30'd758671804;
array[3349]=30'd816348600;
array[3350]=30'd816348600;
array[3351]=30'd798493124;
array[3352]=30'd798493124;
array[3353]=30'd881300969;
array[3354]=30'd916921900;
array[3355]=30'd898043496;
array[3356]=30'd879168118;
array[3357]=30'd879168118;
array[3358]=30'd879168118;
array[3359]=30'd879168118;
array[3360]=30'd898043496;
array[3361]=30'd898043496;
array[3362]=30'd898043496;
array[3363]=30'd898043496;
array[3364]=30'd898043496;
array[3365]=30'd898043496;
array[3366]=30'd959928886;
array[3367]=30'd936883742;
array[3368]=30'd983039487;
array[3369]=30'd983039487;
array[3370]=30'd983039487;
array[3371]=30'd898119130;
array[3372]=30'd798493124;
array[3373]=30'd903304711;
array[3374]=30'd884420162;
array[3375]=30'd898043496;
array[3376]=30'd898043496;
array[3377]=30'd898043496;
array[3378]=30'd842499661;
array[3379]=30'd810005031;
array[3380]=30'd1034407430;
array[3381]=30'd1034407430;
array[3382]=30'd725052963;
array[3383]=30'd938933826;
array[3384]=30'd898043496;
array[3385]=30'd898043496;
array[3386]=30'd898043496;
array[3387]=30'd898043496;
array[3388]=30'd898043496;
array[3389]=30'd898043496;
array[3390]=30'd919054939;
array[3391]=30'd855119431;
array[3392]=30'd827871766;
array[3393]=30'd827871766;
array[3394]=30'd827871766;
array[3395]=30'd857224695;
array[3396]=30'd857224695;
array[3397]=30'd881300969;
array[3398]=30'd960978443;
array[3399]=30'd916921900;
array[3400]=30'd898043496;
array[3401]=30'd879168118;
array[3402]=30'd683036269;
array[3403]=30'd634745492;
array[3404]=30'd608527024;
array[3405]=30'd452327079;
array[3406]=30'd340142721;
array[3407]=30'd289838696;
array[3408]=30'd387329638;
array[3409]=30'd448143984;
array[3410]=30'd408333955;
array[3411]=30'd267838034;
array[3412]=30'd448143984;
array[3413]=30'd448143984;
array[3414]=30'd448143984;
array[3415]=30'd398924382;
array[3416]=30'd259510865;
array[3417]=30'd359106099;
array[3418]=30'd756500033;
array[3419]=30'd815194717;
array[3420]=30'd815194717;
array[3421]=30'd794241637;
array[3422]=30'd709306968;
array[3423]=30'd458750516;
array[3424]=30'd300459585;
array[3425]=30'd300459585;
array[3426]=30'd300459585;
array[3427]=30'd300459585;
array[3428]=30'd323442246;
array[3429]=30'd448143984;
array[3430]=30'd551919254;
array[3431]=30'd427157133;
array[3432]=30'd288811658;
array[3433]=30'd387329638;
array[3434]=30'd361121389;
array[3435]=30'd387329638;
array[3436]=30'd467006094;
array[3437]=30'd551919254;
array[3438]=30'd729186945;
array[3439]=30'd898043496;
array[3440]=30'd898043496;
array[3441]=30'd898043496;
array[3442]=30'd919054939;
array[3443]=30'd877139478;
array[3444]=30'd785935846;
array[3445]=30'd798493124;
array[3446]=30'd798493124;
array[3447]=30'd821544417;
array[3448]=30'd821544417;
array[3449]=30'd860309028;
array[3450]=30'd884420162;
array[3451]=30'd879168118;
array[3452]=30'd898043496;
array[3453]=30'd879168118;
array[3454]=30'd879168118;
array[3455]=30'd879168118;
array[3456]=30'd898043496;
array[3457]=30'd898043496;
array[3458]=30'd898043496;
array[3459]=30'd898043496;
array[3460]=30'd898043496;
array[3461]=30'd919054939;
array[3462]=30'd936883742;
array[3463]=30'd877139478;
array[3464]=30'd857224695;
array[3465]=30'd903304711;
array[3466]=30'd921177592;
array[3467]=30'd1016593896;
array[3468]=30'd871910847;
array[3469]=30'd821544417;
array[3470]=30'd903304711;
array[3471]=30'd938933826;
array[3472]=30'd898043496;
array[3473]=30'd898043496;
array[3474]=30'd898043496;
array[3475]=30'd779606588;
array[3476]=30'd1034407430;
array[3477]=30'd1034407430;
array[3478]=30'd810005031;
array[3479]=30'd884420162;
array[3480]=30'd898043496;
array[3481]=30'd898043496;
array[3482]=30'd898043496;
array[3483]=30'd898043496;
array[3484]=30'd898043496;
array[3485]=30'd919054939;
array[3486]=30'd855119431;
array[3487]=30'd827871766;
array[3488]=30'd921177592;
array[3489]=30'd964180446;
array[3490]=30'd921177592;
array[3491]=30'd898119130;
array[3492]=30'd833115609;
array[3493]=30'd881300969;
array[3494]=30'd945268200;
array[3495]=30'd916921900;
array[3496]=30'd898043496;
array[3497]=30'd879168118;
array[3498]=30'd624350812;
array[3499]=30'd634745492;
array[3500]=30'd613805729;
array[3501]=30'd427157133;
array[3502]=30'd340142721;
array[3503]=30'd318144090;
array[3504]=30'd361121389;
array[3505]=30'd448143984;
array[3506]=30'd408333955;
array[3507]=30'd239530594;
array[3508]=30'd448143984;
array[3509]=30'd448143984;
array[3510]=30'd398924382;
array[3511]=30'd302486106;
array[3512]=30'd300459585;
array[3513]=30'd354967120;
array[3514]=30'd694642226;
array[3515]=30'd815194717;
array[3516]=30'd794241637;
array[3517]=30'd592910950;
array[3518]=30'd283619908;
array[3519]=30'd300459585;
array[3520]=30'd282664514;
array[3521]=30'd282664514;
array[3522]=30'd282664514;
array[3523]=30'd300459585;
array[3524]=30'd341225034;
array[3525]=30'd558250630;
array[3526]=30'd467006094;
array[3527]=30'd408333955;
array[3528]=30'd289838696;
array[3529]=30'd408333955;
array[3530]=30'd318144090;
array[3531]=30'd387329638;
array[3532]=30'd467006094;
array[3533]=30'd522581659;
array[3534]=30'd781608573;
array[3535]=30'd898043496;
array[3536]=30'd898043496;
array[3537]=30'd898043496;
array[3538]=30'd898043496;
array[3539]=30'd919054939;
array[3540]=30'd898098744;
array[3541]=30'd884420162;
array[3542]=30'd860309028;
array[3543]=30'd916921900;
array[3544]=30'd884420162;
array[3545]=30'd898043496;
array[3546]=30'd898043496;
array[3547]=30'd898043496;
array[3548]=30'd898043496;
array[3549]=30'd879168118;
array[3550]=30'd879168118;
array[3551]=30'd898043496;
array[3552]=30'd898043496;
array[3553]=30'd898043496;
array[3554]=30'd898043496;
array[3555]=30'd898043496;
array[3556]=30'd919054939;
array[3557]=30'd898098744;
array[3558]=30'd827871766;
array[3559]=30'd785935846;
array[3560]=30'd798493124;
array[3561]=30'd798493124;
array[3562]=30'd821544417;
array[3563]=30'd964180446;
array[3564]=30'd983039487;
array[3565]=30'd833115609;
array[3566]=30'd821544417;
array[3567]=30'd916921900;
array[3568]=30'd919054939;
array[3569]=30'd884420162;
array[3570]=30'd842499661;
array[3571]=30'd725052963;
array[3572]=30'd1034407430;
array[3573]=30'd1034407430;
array[3574]=30'd903304711;
array[3575]=30'd795279924;
array[3576]=30'd898043496;
array[3577]=30'd898043496;
array[3578]=30'd898043496;
array[3579]=30'd898043496;
array[3580]=30'd919054939;
array[3581]=30'd877139478;
array[3582]=30'd827871766;
array[3583]=30'd964180446;
array[3584]=30'd983039487;
array[3585]=30'd921177592;
array[3586]=30'd898119130;
array[3587]=30'd898119130;
array[3588]=30'd898119130;
array[3589]=30'd852996553;
array[3590]=30'd945268200;
array[3591]=30'd916921900;
array[3592]=30'd898043496;
array[3593]=30'd898043496;
array[3594]=30'd624350812;
array[3595]=30'd634745492;
array[3596]=30'd559255224;
array[3597]=30'd393597595;
array[3598]=30'd340142721;
array[3599]=30'd361121389;
array[3600]=30'd344392301;
array[3601]=30'd448143984;
array[3602]=30'd459725411;
array[3603]=30'd341225034;
array[3604]=30'd344392301;
array[3605]=30'd341225034;
array[3606]=30'd283619908;
array[3607]=30'd300459585;
array[3608]=30'd300459585;
array[3609]=30'd354967120;
array[3610]=30'd779606588;
array[3611]=30'd756500033;
array[3612]=30'd506974798;
array[3613]=30'd259510865;
array[3614]=30'd300459585;
array[3615]=30'd282664514;
array[3616]=30'd282664514;
array[3617]=30'd282664514;
array[3618]=30'd300459585;
array[3619]=30'd259510865;
array[3620]=30'd448143984;
array[3621]=30'd522581659;
array[3622]=30'd393597595;
array[3623]=30'd289838696;
array[3624]=30'd344392301;
array[3625]=30'd459725411;
array[3626]=30'd318144090;
array[3627]=30'd387329638;
array[3628]=30'd467006094;
array[3629]=30'd522581659;
array[3630]=30'd815194717;
array[3631]=30'd898043496;
array[3632]=30'd898043496;
array[3633]=30'd898043496;
array[3634]=30'd898043496;
array[3635]=30'd898043496;
array[3636]=30'd898043496;
array[3637]=30'd898043496;
array[3638]=30'd898043496;
array[3639]=30'd898043496;
array[3640]=30'd898043496;
array[3641]=30'd898043496;
array[3642]=30'd898043496;
array[3643]=30'd898043496;
array[3644]=30'd879168118;
array[3645]=30'd879168118;
array[3646]=30'd879168118;
array[3647]=30'd898043496;
array[3648]=30'd898043496;
array[3649]=30'd898043496;
array[3650]=30'd898043496;
array[3651]=30'd898043496;
array[3652]=30'd919054939;
array[3653]=30'd936883742;
array[3654]=30'd833115609;
array[3655]=30'd945316283;
array[3656]=30'd945316283;
array[3657]=30'd911766951;
array[3658]=30'd798493124;
array[3659]=30'd881300969;
array[3660]=30'd983039487;
array[3661]=30'd925360587;
array[3662]=30'd798493124;
array[3663]=30'd903304711;
array[3664]=30'd936883742;
array[3665]=30'd827871766;
array[3666]=30'd821544417;
array[3667]=30'd693598700;
array[3668]=30'd1034407430;
array[3669]=30'd1034407430;
array[3670]=30'd936883742;
array[3671]=30'd756500033;
array[3672]=30'd919054939;
array[3673]=30'd898043496;
array[3674]=30'd898043496;
array[3675]=30'd898043496;
array[3676]=30'd898098744;
array[3677]=30'd827871766;
array[3678]=30'd964180446;
array[3679]=30'd964180446;
array[3680]=30'd857224695;
array[3681]=30'd833115609;
array[3682]=30'd833115609;
array[3683]=30'd833115609;
array[3684]=30'd871910847;
array[3685]=30'd871910847;
array[3686]=30'd881300969;
array[3687]=30'd916921900;
array[3688]=30'd884420162;
array[3689]=30'd898043496;
array[3690]=30'd592910950;
array[3691]=30'd634745492;
array[3692]=30'd551919254;
array[3693]=30'd340142721;
array[3694]=30'd289838696;
array[3695]=30'd414594647;
array[3696]=30'd344392301;
array[3697]=30'd344392301;
array[3698]=30'd344392301;
array[3699]=30'd259510865;
array[3700]=30'd259510865;
array[3701]=30'd236450390;
array[3702]=30'd300459585;
array[3703]=30'd300459585;
array[3704]=30'd282664514;
array[3705]=30'd335057455;
array[3706]=30'd725091917;
array[3707]=30'd444087878;
array[3708]=30'd252253768;
array[3709]=30'd300459585;
array[3710]=30'd282664514;
array[3711]=30'd282664514;
array[3712]=30'd282664514;
array[3713]=30'd282664514;
array[3714]=30'd300459585;
array[3715]=30'd259510865;
array[3716]=30'd558250630;
array[3717]=30'd467006094;
array[3718]=30'd387329638;
array[3719]=30'd239530594;
array[3720]=30'd289838696;
array[3721]=30'd344392301;
array[3722]=30'd289838696;
array[3723]=30'd387329638;
array[3724]=30'd485876339;
array[3725]=30'd522581659;
array[3726]=30'd815194717;
array[3727]=30'd898043496;
array[3728]=30'd898043496;
array[3729]=30'd898043496;
array[3730]=30'd898043496;
array[3731]=30'd879168118;
array[3732]=30'd898043496;
array[3733]=30'd879168118;
array[3734]=30'd898043496;
array[3735]=30'd898043496;
array[3736]=30'd898043496;
array[3737]=30'd879168118;
array[3738]=30'd879168118;
array[3739]=30'd898043496;
array[3740]=30'd898043496;
array[3741]=30'd898043496;
array[3742]=30'd879168118;
array[3743]=30'd898043496;
array[3744]=30'd898043496;
array[3745]=30'd898043496;
array[3746]=30'd898043496;
array[3747]=30'd919054939;
array[3748]=30'd898098744;
array[3749]=30'd877139478;
array[3750]=30'd816348600;
array[3751]=30'd850952611;
array[3752]=30'd850952611;
array[3753]=30'd945316283;
array[3754]=30'd816348600;
array[3755]=30'd852996553;
array[3756]=30'd921177592;
array[3757]=30'd898119130;
array[3758]=30'd798493124;
array[3759]=30'd903304711;
array[3760]=30'd936883742;
array[3761]=30'd983039487;
array[3762]=30'd983039487;
array[3763]=30'd706223587;
array[3764]=30'd1000848926;
array[3765]=30'd1034407430;
array[3766]=30'd1000848926;
array[3767]=30'd725052963;
array[3768]=30'd919054939;
array[3769]=30'd898043496;
array[3770]=30'd898043496;
array[3771]=30'd919054939;
array[3772]=30'd855119431;
array[3773]=30'd857224695;
array[3774]=30'd964180446;
array[3775]=30'd857224695;
array[3776]=30'd833115609;
array[3777]=30'd898119130;
array[3778]=30'd945316283;
array[3779]=30'd945316283;
array[3780]=30'd816348600;
array[3781]=30'd911766951;
array[3782]=30'd852996553;
array[3783]=30'd960978443;
array[3784]=30'd884420162;
array[3785]=30'd898043496;
array[3786]=30'd566698607;
array[3787]=30'd634745492;
array[3788]=30'd551919254;
array[3789]=30'd340142721;
array[3790]=30'd289838696;
array[3791]=30'd344392301;
array[3792]=30'd391685709;
array[3793]=30'd452485730;
array[3794]=30'd482898518;
array[3795]=30'd314134080;
array[3796]=30'd282664514;
array[3797]=30'd244888116;
array[3798]=30'd282664514;
array[3799]=30'd282664514;
array[3800]=30'd282664514;
array[3801]=30'd252253768;
array[3802]=30'd335057455;
array[3803]=30'd300459585;
array[3804]=30'd300459585;
array[3805]=30'd282664514;
array[3806]=30'd282664514;
array[3807]=30'd282664514;
array[3808]=30'd282664514;
array[3809]=30'd282664514;
array[3810]=30'd244888116;
array[3811]=30'd459725411;
array[3812]=30'd527847013;
array[3813]=30'd427157133;
array[3814]=30'd288811658;
array[3815]=30'd239530594;
array[3816]=30'd283619908;
array[3817]=30'd259510865;
array[3818]=30'd230137397;
array[3819]=30'd341225034;
array[3820]=30'd448143984;
array[3821]=30'd527847013;
array[3822]=30'd794241637;
array[3823]=30'd898043496;
array[3824]=30'd898043496;
array[3825]=30'd898043496;
array[3826]=30'd898043496;
array[3827]=30'd898043496;
array[3828]=30'd898043496;
array[3829]=30'd898043496;
array[3830]=30'd898043496;
array[3831]=30'd898043496;
array[3832]=30'd898043496;
array[3833]=30'd898043496;
array[3834]=30'd879168118;
array[3835]=30'd898043496;
array[3836]=30'd898043496;
array[3837]=30'd898043496;
array[3838]=30'd898043496;
array[3839]=30'd898043496;
array[3840]=30'd898043496;
array[3841]=30'd898043496;
array[3842]=30'd898043496;
array[3843]=30'd919054939;
array[3844]=30'd936883742;
array[3845]=30'd833115609;
array[3846]=30'd850952611;
array[3847]=30'd790145435;
array[3848]=30'd816348600;
array[3849]=30'd911766951;
array[3850]=30'd816348600;
array[3851]=30'd852996553;
array[3852]=30'd921177592;
array[3853]=30'd898119130;
array[3854]=30'd798493124;
array[3855]=30'd903304711;
array[3856]=30'd877139478;
array[3857]=30'd857224695;
array[3858]=30'd898119130;
array[3859]=30'd706223587;
array[3860]=30'd983039487;
array[3861]=30'd1034407430;
array[3862]=30'd1034407430;
array[3863]=30'd725052963;
array[3864]=30'd938933826;
array[3865]=30'd919054939;
array[3866]=30'd919054939;
array[3867]=30'd919054939;
array[3868]=30'd877139478;
array[3869]=30'd857224695;
array[3870]=30'd964180446;
array[3871]=30'd833115609;
array[3872]=30'd898119130;
array[3873]=30'd945316283;
array[3874]=30'd816348600;
array[3875]=30'd850952611;
array[3876]=30'd790145435;
array[3877]=30'd911766951;
array[3878]=30'd816348600;
array[3879]=30'd960978443;
array[3880]=30'd884420162;
array[3881]=30'd898043496;
array[3882]=30'd527847013;
array[3883]=30'd634745492;
array[3884]=30'd522581659;
array[3885]=30'd288811658;
array[3886]=30'd354967120;
array[3887]=30'd482898518;
array[3888]=30'd473528913;
array[3889]=30'd473528913;
array[3890]=30'd473528913;
array[3891]=30'd370760263;
array[3892]=30'd282664514;
array[3893]=30'd252253768;
array[3894]=30'd282664514;
array[3895]=30'd282664514;
array[3896]=30'd282664514;
array[3897]=30'd252253768;
array[3898]=30'd252253768;
array[3899]=30'd300459585;
array[3900]=30'd282664514;
array[3901]=30'd282664514;
array[3902]=30'd282664514;
array[3903]=30'd314134080;
array[3904]=30'd282664514;
array[3905]=30'd300459585;
array[3906]=30'd323442246;
array[3907]=30'd559303250;
array[3908]=30'd427157133;
array[3909]=30'd408333955;
array[3910]=30'd289838696;
array[3911]=30'd302486106;
array[3912]=30'd354967120;
array[3913]=30'd346647116;
array[3914]=30'd391685709;
array[3915]=30'd354967120;
array[3916]=30'd377963103;
array[3917]=30'd527847013;
array[3918]=30'd729186945;
array[3919]=30'd898043496;
array[3920]=30'd898043496;
array[3921]=30'd898043496;
array[3922]=30'd898043496;
array[3923]=30'd898043496;
array[3924]=30'd898043496;
array[3925]=30'd898043496;
array[3926]=30'd898043496;
array[3927]=30'd898043496;
array[3928]=30'd898043496;
array[3929]=30'd898043496;
array[3930]=30'd898043496;
array[3931]=30'd898043496;
array[3932]=30'd898043496;
array[3933]=30'd898043496;
array[3934]=30'd898043496;
array[3935]=30'd879168118;
array[3936]=30'd898043496;
array[3937]=30'd919054939;
array[3938]=30'd898043496;
array[3939]=30'd919054939;
array[3940]=30'd936883742;
array[3941]=30'd833115609;
array[3942]=30'd885566856;
array[3943]=30'd850952611;
array[3944]=30'd850952611;
array[3945]=30'd949526930;
array[3946]=30'd871910847;
array[3947]=30'd798493124;
array[3948]=30'd921177592;
array[3949]=30'd898119130;
array[3950]=30'd821544417;
array[3951]=30'd945268200;
array[3952]=30'd821544417;
array[3953]=30'd758671804;
array[3954]=30'd740803022;
array[3955]=30'd621275606;
array[3956]=30'd821544417;
array[3957]=30'd843548160;
array[3958]=30'd746067471;
array[3959]=30'd555187752;
array[3960]=30'd810005031;
array[3961]=30'd842499661;
array[3962]=30'd799523423;
array[3963]=30'd898098744;
array[3964]=30'd898098744;
array[3965]=30'd827871766;
array[3966]=30'd921177592;
array[3967]=30'd857224695;
array[3968]=30'd857224695;
array[3969]=30'd898119130;
array[3970]=30'd816348600;
array[3971]=30'd850952611;
array[3972]=30'd850952611;
array[3973]=30'd816348600;
array[3974]=30'd881300969;
array[3975]=30'd960978443;
array[3976]=30'd884420162;
array[3977]=30'd898043496;
array[3978]=30'd566698607;
array[3979]=30'd634745492;
array[3980]=30'd496374434;
array[3981]=30'd289838696;
array[3982]=30'd421031501;
array[3983]=30'd461984322;
array[3984]=30'd488205898;
array[3985]=30'd473528913;
array[3986]=30'd473528913;
array[3987]=30'd461984322;
array[3988]=30'd314134080;
array[3989]=30'd252253768;
array[3990]=30'd282664514;
array[3991]=30'd282664514;
array[3992]=30'd282664514;
array[3993]=30'd220784191;
array[3994]=30'd220784191;
array[3995]=30'd282664514;
array[3996]=30'd282664514;
array[3997]=30'd282664514;
array[3998]=30'd282664514;
array[3999]=30'd282664514;
array[4000]=30'd282664514;
array[4001]=30'd244888116;
array[4002]=30'd459725411;
array[4003]=30'd483822211;
array[4004]=30'd427157133;
array[4005]=30'd344392301;
array[4006]=30'd344392301;
array[4007]=30'd444087878;
array[4008]=30'd461984322;
array[4009]=30'd461984322;
array[4010]=30'd461984322;
array[4011]=30'd478743092;
array[4012]=30'd421031501;
array[4013]=30'd398924382;
array[4014]=30'd709306968;
array[4015]=30'd898043496;
array[4016]=30'd898043496;
array[4017]=30'd898043496;
array[4018]=30'd898043496;
array[4019]=30'd898043496;
array[4020]=30'd898043496;
array[4021]=30'd898043496;
array[4022]=30'd898043496;
array[4023]=30'd898043496;
array[4024]=30'd898043496;
array[4025]=30'd898043496;
array[4026]=30'd898043496;
array[4027]=30'd898043496;
array[4028]=30'd898043496;
array[4029]=30'd898043496;
array[4030]=30'd898043496;
array[4031]=30'd898043496;
array[4032]=30'd898043496;
array[4033]=30'd898043496;
array[4034]=30'd919054939;
array[4035]=30'd919054939;
array[4036]=30'd959928886;
array[4037]=30'd898119130;
array[4038]=30'd816348600;
array[4039]=30'd850952611;
array[4040]=30'd774396326;
array[4041]=30'd790145435;
array[4042]=30'd816348600;
array[4043]=30'd871910847;
array[4044]=30'd925360587;
array[4045]=30'd833115609;
array[4046]=30'd881300969;
array[4047]=30'd945268200;
array[4048]=30'd921177592;
array[4049]=30'd706223587;
array[4050]=30'd649571855;
array[4051]=30'd770126332;
array[4052]=30'd903304711;
array[4053]=30'd936883742;
array[4054]=30'd936883742;
array[4055]=30'd916921900;
array[4056]=30'd810005031;
array[4057]=30'd612873765;
array[4058]=30'd810005031;
array[4059]=30'd668430907;
array[4060]=30'd898098744;
array[4061]=30'd877139478;
array[4062]=30'd936883742;
array[4063]=30'd921177592;
array[4064]=30'd857224695;
array[4065]=30'd833115609;
array[4066]=30'd816348600;
array[4067]=30'd850952611;
array[4068]=30'd850952611;
array[4069]=30'd945316283;
array[4070]=30'd945268200;
array[4071]=30'd916921900;
array[4072]=30'd898043496;
array[4073]=30'd898043496;
array[4074]=30'd592910950;
array[4075]=30'd653676161;
array[4076]=30'd483822211;
array[4077]=30'd302486106;
array[4078]=30'd452485730;
array[4079]=30'd461984322;
array[4080]=30'd488205898;
array[4081]=30'd473528913;
array[4082]=30'd488205898;
array[4083]=30'd473528913;
array[4084]=30'd346647116;
array[4085]=30'd282664514;
array[4086]=30'd282664514;
array[4087]=30'd282664514;
array[4088]=30'd220784191;
array[4089]=30'd252253768;
array[4090]=30'd220784191;
array[4091]=30'd252253768;
array[4092]=30'd282664514;
array[4093]=30'd282664514;
array[4094]=30'd282664514;
array[4095]=30'd282664514;
array[4096]=30'd282664514;
array[4097]=30'd283619908;
array[4098]=30'd527847013;
array[4099]=30'd434534016;
array[4100]=30'd387329638;
array[4101]=30'd344392301;
array[4102]=30'd377963103;
array[4103]=30'd482898518;
array[4104]=30'd461984322;
array[4105]=30'd473528913;
array[4106]=30'd473528913;
array[4107]=30'd473528913;
array[4108]=30'd461984322;
array[4109]=30'd421031501;
array[4110]=30'd612873765;
array[4111]=30'd919054939;
array[4112]=30'd898043496;
array[4113]=30'd898043496;
array[4114]=30'd898043496;
array[4115]=30'd898043496;
array[4116]=30'd898043496;
array[4117]=30'd898043496;
array[4118]=30'd898043496;
array[4119]=30'd898043496;
array[4120]=30'd898043496;
array[4121]=30'd898043496;
array[4122]=30'd898043496;
array[4123]=30'd898043496;
array[4124]=30'd898043496;
array[4125]=30'd898043496;
array[4126]=30'd898043496;
array[4127]=30'd898043496;
array[4128]=30'd898043496;
array[4129]=30'd898043496;
array[4130]=30'd919054939;
array[4131]=30'd919054939;
array[4132]=30'd959928886;
array[4133]=30'd983039487;
array[4134]=30'd816348600;
array[4135]=30'd832088453;
array[4136]=30'd850952611;
array[4137]=30'd911766951;
array[4138]=30'd911766951;
array[4139]=30'd871910847;
array[4140]=30'd833115609;
array[4141]=30'd833115609;
array[4142]=30'd857224695;
array[4143]=30'd857224695;
array[4144]=30'd821544417;
array[4145]=30'd843548160;
array[4146]=30'd960978443;
array[4147]=30'd959928886;
array[4148]=30'd979842606;
array[4149]=30'd979842606;
array[4150]=30'd959928886;
array[4151]=30'd959928886;
array[4152]=30'd936883742;
array[4153]=30'd756500033;
array[4154]=30'd979842606;
array[4155]=30'd725052963;
array[4156]=30'd898098744;
array[4157]=30'd959928886;
array[4158]=30'd898098744;
array[4159]=30'd898098744;
array[4160]=30'd898098744;
array[4161]=30'd936883742;
array[4162]=30'd921177592;
array[4163]=30'd921177592;
array[4164]=30'd983039487;
array[4165]=30'd960978443;
array[4166]=30'd916921900;
array[4167]=30'd898043496;
array[4168]=30'd898043496;
array[4169]=30'd898043496;
array[4170]=30'd548890196;
array[4171]=30'd625322602;
array[4172]=30'd483822211;
array[4173]=30'd302486106;
array[4174]=30'd482898518;
array[4175]=30'd473528913;
array[4176]=30'd473528913;
array[4177]=30'd488205898;
array[4178]=30'd473528913;
array[4179]=30'd473528913;
array[4180]=30'd370760263;
array[4181]=30'd282664514;
array[4182]=30'd252253768;
array[4183]=30'd252253768;
array[4184]=30'd198780482;
array[4185]=30'd220784191;
array[4186]=30'd244888116;
array[4187]=30'd244888116;
array[4188]=30'd252253768;
array[4189]=30'd282664514;
array[4190]=30'd282664514;
array[4191]=30'd314134080;
array[4192]=30'd370760263;
array[4193]=30'd359106099;
array[4194]=30'd558250630;
array[4195]=30'd408333955;
array[4196]=30'd267838034;
array[4197]=30'd398924382;
array[4198]=30'd354967120;
array[4199]=30'd482898518;
array[4200]=30'd473528913;
array[4201]=30'd473528913;
array[4202]=30'd473528913;
array[4203]=30'd461984322;
array[4204]=30'd434727495;
array[4205]=30'd434727495;
array[4206]=30'd444087878;
array[4207]=30'd799523423;
array[4208]=30'd898043496;
array[4209]=30'd898043496;
array[4210]=30'd898043496;
array[4211]=30'd919054939;
array[4212]=30'd898043496;
array[4213]=30'd898043496;
array[4214]=30'd898043496;
array[4215]=30'd898043496;
array[4216]=30'd898043496;
array[4217]=30'd898043496;
array[4218]=30'd898043496;
array[4219]=30'd898043496;
array[4220]=30'd898043496;
array[4221]=30'd898043496;
array[4222]=30'd898043496;
array[4223]=30'd898043496;
array[4224]=30'd898043496;
array[4225]=30'd898043496;
array[4226]=30'd919054939;
array[4227]=30'd919054939;
array[4228]=30'd919054939;
array[4229]=30'd1000848926;
array[4230]=30'd898119130;
array[4231]=30'd790145435;
array[4232]=30'd850952611;
array[4233]=30'd816348600;
array[4234]=30'd790145435;
array[4235]=30'd816348600;
array[4236]=30'd871910847;
array[4237]=30'd921177592;
array[4238]=30'd898119130;
array[4239]=30'd775423471;
array[4240]=30'd621275606;
array[4241]=30'd945268200;
array[4242]=30'd960978443;
array[4243]=30'd959928886;
array[4244]=30'd959928886;
array[4245]=30'd979842606;
array[4246]=30'd979842606;
array[4247]=30'd959928886;
array[4248]=30'd936883742;
array[4249]=30'd725052963;
array[4250]=30'd979842606;
array[4251]=30'd725052963;
array[4252]=30'd938933826;
array[4253]=30'd919054939;
array[4254]=30'd919054939;
array[4255]=30'd919054939;
array[4256]=30'd919054939;
array[4257]=30'd919054939;
array[4258]=30'd919054939;
array[4259]=30'd898098744;
array[4260]=30'd959928886;
array[4261]=30'd938933826;
array[4262]=30'd938933826;
array[4263]=30'd898043496;
array[4264]=30'd898043496;
array[4265]=30'd799523423;
array[4266]=30'd377963103;
array[4267]=30'd559303250;
array[4268]=30'd496412259;
array[4269]=30'd302486106;
array[4270]=30'd482898518;
array[4271]=30'd488205898;
array[4272]=30'd488205898;
array[4273]=30'd488205898;
array[4274]=30'd473528913;
array[4275]=30'd473528913;
array[4276]=30'd434727495;
array[4277]=30'd314134080;
array[4278]=30'd314134080;
array[4279]=30'd282664514;
array[4280]=30'd252253768;
array[4281]=30'd220784191;
array[4282]=30'd282664514;
array[4283]=30'd314134080;
array[4284]=30'd282664514;
array[4285]=30'd370760263;
array[4286]=30'd434727495;
array[4287]=30'd434727495;
array[4288]=30'd314134080;
array[4289]=30'd428280389;
array[4290]=30'd527847013;
array[4291]=30'd398924382;
array[4292]=30'd213323368;
array[4293]=30'd377963103;
array[4294]=30'd391685709;
array[4295]=30'd482898518;
array[4296]=30'd473528913;
array[4297]=30'd473528913;
array[4298]=30'd473528913;
array[4299]=30'd434727495;
array[4300]=30'd370760263;
array[4301]=30'd473528913;
array[4302]=30'd478743092;
array[4303]=30'd562592331;
array[4304]=30'd919054939;
array[4305]=30'd919054939;
array[4306]=30'd898043496;
array[4307]=30'd898043496;
array[4308]=30'd898043496;
array[4309]=30'd898043496;
array[4310]=30'd898043496;
array[4311]=30'd898043496;
array[4312]=30'd898043496;
array[4313]=30'd898043496;
array[4314]=30'd898043496;
array[4315]=30'd898043496;
array[4316]=30'd898043496;
array[4317]=30'd898043496;
array[4318]=30'd898043496;
array[4319]=30'd898043496;
array[4320]=30'd919054939;
array[4321]=30'd919054939;
array[4322]=30'd919054939;
array[4323]=30'd919054939;
array[4324]=30'd919054939;
array[4325]=30'd959928886;
array[4326]=30'd983039487;
array[4327]=30'd921177592;
array[4328]=30'd871910847;
array[4329]=30'd871910847;
array[4330]=30'd925360587;
array[4331]=30'd964180446;
array[4332]=30'd921177592;
array[4333]=30'd936883742;
array[4334]=30'd983039487;
array[4335]=30'd921177592;
array[4336]=30'd596111858;
array[4337]=30'd960978443;
array[4338]=30'd960978443;
array[4339]=30'd959928886;
array[4340]=30'd959928886;
array[4341]=30'd979842606;
array[4342]=30'd979842606;
array[4343]=30'd959928886;
array[4344]=30'd959928886;
array[4345]=30'd795279924;
array[4346]=30'd936883742;
array[4347]=30'd694642226;
array[4348]=30'd919054939;
array[4349]=30'd919054939;
array[4350]=30'd919054939;
array[4351]=30'd919054939;
array[4352]=30'd919054939;
array[4353]=30'd919054939;
array[4354]=30'd919054939;
array[4355]=30'd919054939;
array[4356]=30'd919054939;
array[4357]=30'd938933826;
array[4358]=30'd898043496;
array[4359]=30'd919054939;
array[4360]=30'd898043496;
array[4361]=30'd562592331;
array[4362]=30'd444087878;
array[4363]=30'd459725411;
array[4364]=30'd496412259;
array[4365]=30'd359106099;
array[4366]=30'd482898518;
array[4367]=30'd488205898;
array[4368]=30'd488205898;
array[4369]=30'd488205898;
array[4370]=30'd473528913;
array[4371]=30'd473528913;
array[4372]=30'd473528913;
array[4373]=30'd473528913;
array[4374]=30'd461984322;
array[4375]=30'd461984322;
array[4376]=30'd370760263;
array[4377]=30'd282664514;
array[4378]=30'd434727495;
array[4379]=30'd461984322;
array[4380]=30'd461984322;
array[4381]=30'd370760263;
array[4382]=30'd370760263;
array[4383]=30'd370760263;
array[4384]=30'd421031501;
array[4385]=30'd475488805;
array[4386]=30'd459725411;
array[4387]=30'd289838696;
array[4388]=30'd236450390;
array[4389]=30'd354967120;
array[4390]=30'd444087878;
array[4391]=30'd461984322;
array[4392]=30'd473528913;
array[4393]=30'd473528913;
array[4394]=30'd461984322;
array[4395]=30'd370760263;
array[4396]=30'd461984322;
array[4397]=30'd473528913;
array[4398]=30'd473528913;
array[4399]=30'd434727495;
array[4400]=30'd842499661;
array[4401]=30'd919054939;
array[4402]=30'd898043496;
array[4403]=30'd898043496;
array[4404]=30'd898043496;
array[4405]=30'd898043496;
array[4406]=30'd898043496;
array[4407]=30'd898043496;
array[4408]=30'd898043496;
array[4409]=30'd898043496;
array[4410]=30'd898043496;
array[4411]=30'd898043496;
array[4412]=30'd898043496;
array[4413]=30'd898043496;
array[4414]=30'd898043496;
array[4415]=30'd898043496;
array[4416]=30'd919054939;
array[4417]=30'd919054939;
array[4418]=30'd919054939;
array[4419]=30'd919054939;
array[4420]=30'd919054939;
array[4421]=30'd919054939;
array[4422]=30'd919054939;
array[4423]=30'd959928886;
array[4424]=30'd936883742;
array[4425]=30'd936883742;
array[4426]=30'd936883742;
array[4427]=30'd936883742;
array[4428]=30'd898098744;
array[4429]=30'd898098744;
array[4430]=30'd919054939;
array[4431]=30'd1000848926;
array[4432]=30'd725052963;
array[4433]=30'd936883742;
array[4434]=30'd959928886;
array[4435]=30'd959928886;
array[4436]=30'd959928886;
array[4437]=30'd979842606;
array[4438]=30'd979842606;
array[4439]=30'd959928886;
array[4440]=30'd959928886;
array[4441]=30'd916921900;
array[4442]=30'd612873765;
array[4443]=30'd884420162;
array[4444]=30'd919054939;
array[4445]=30'd919054939;
array[4446]=30'd919054939;
array[4447]=30'd919054939;
array[4448]=30'd919054939;
array[4449]=30'd919054939;
array[4450]=30'd919054939;
array[4451]=30'd919054939;
array[4452]=30'd919054939;
array[4453]=30'd919054939;
array[4454]=30'd919054939;
array[4455]=30'd919054939;
array[4456]=30'd799523423;
array[4457]=30'd444087878;
array[4458]=30'd482898518;
array[4459]=30'd354967120;
array[4460]=30'd506974798;
array[4461]=30'd332951128;
array[4462]=30'd482898518;
array[4463]=30'd461984322;
array[4464]=30'd488205898;
array[4465]=30'd488205898;
array[4466]=30'd488205898;
array[4467]=30'd488205898;
array[4468]=30'd488205898;
array[4469]=30'd473528913;
array[4470]=30'd473528913;
array[4471]=30'd473528913;
array[4472]=30'd434727495;
array[4473]=30'd370760263;
array[4474]=30'd473528913;
array[4475]=30'd473528913;
array[4476]=30'd473528913;
array[4477]=30'd473528913;
array[4478]=30'd461984322;
array[4479]=30'd461984322;
array[4480]=30'd478743092;
array[4481]=30'd458750516;
array[4482]=30'd398924382;
array[4483]=30'd302486106;
array[4484]=30'd391685709;
array[4485]=30'd300459585;
array[4486]=30'd421031501;
array[4487]=30'd473528913;
array[4488]=30'd473528913;
array[4489]=30'd473528913;
array[4490]=30'd434727495;
array[4491]=30'd434727495;
array[4492]=30'd473528913;
array[4493]=30'd473528913;
array[4494]=30'd473528913;
array[4495]=30'd461984322;
array[4496]=30'd725091917;
array[4497]=30'd919054939;
array[4498]=30'd898043496;
array[4499]=30'd898043496;
array[4500]=30'd898043496;
array[4501]=30'd898043496;
array[4502]=30'd898043496;
array[4503]=30'd898043496;
array[4504]=30'd898043496;
array[4505]=30'd898043496;
array[4506]=30'd898043496;
array[4507]=30'd898043496;
array[4508]=30'd898043496;
array[4509]=30'd898043496;
array[4510]=30'd898043496;
array[4511]=30'd919054939;
array[4512]=30'd919054939;
array[4513]=30'd919054939;
array[4514]=30'd919054939;
array[4515]=30'd919054939;
array[4516]=30'd919054939;
array[4517]=30'd919054939;
array[4518]=30'd919054939;
array[4519]=30'd919054939;
array[4520]=30'd919054939;
array[4521]=30'd919054939;
array[4522]=30'd919054939;
array[4523]=30'd919054939;
array[4524]=30'd919054939;
array[4525]=30'd919054939;
array[4526]=30'd919054939;
array[4527]=30'd959928886;
array[4528]=30'd810005031;
array[4529]=30'd884420162;
array[4530]=30'd979842606;
array[4531]=30'd979842606;
array[4532]=30'd979842606;
array[4533]=30'd979842606;
array[4534]=30'd979842606;
array[4535]=30'd959928886;
array[4536]=30'd959928886;
array[4537]=30'd959928886;
array[4538]=30'd795279924;
array[4539]=30'd938933826;
array[4540]=30'd919054939;
array[4541]=30'd919054939;
array[4542]=30'd919054939;
array[4543]=30'd919054939;
array[4544]=30'd919054939;
array[4545]=30'd919054939;
array[4546]=30'd919054939;
array[4547]=30'd919054939;
array[4548]=30'd919054939;
array[4549]=30'd919054939;
array[4550]=30'd919054939;
array[4551]=30'd898098744;
array[4552]=30'd482898518;
array[4553]=30'd461984322;
array[4554]=30'd473528913;
array[4555]=30'd482898518;
array[4556]=30'd354967120;
array[4557]=30'd332951128;
array[4558]=30'd391685709;
array[4559]=30'd461984322;
array[4560]=30'd488205898;
array[4561]=30'd488205898;
array[4562]=30'd488205898;
array[4563]=30'd488205898;
array[4564]=30'd488205898;
array[4565]=30'd473528913;
array[4566]=30'd473528913;
array[4567]=30'd473528913;
array[4568]=30'd370760263;
array[4569]=30'd461984322;
array[4570]=30'd473528913;
array[4571]=30'd488205898;
array[4572]=30'd488205898;
array[4573]=30'd488205898;
array[4574]=30'd473528913;
array[4575]=30'd473528913;
array[4576]=30'd461984322;
array[4577]=30'd332951128;
array[4578]=30'd354967120;
array[4579]=30'd391685709;
array[4580]=30'd482898518;
array[4581]=30'd373855782;
array[4582]=30'd370760263;
array[4583]=30'd473528913;
array[4584]=30'd473528913;
array[4585]=30'd461984322;
array[4586]=30'd370760263;
array[4587]=30'd473528913;
array[4588]=30'd473528913;
array[4589]=30'd473528913;
array[4590]=30'd473528913;
array[4591]=30'd461984322;
array[4592]=30'd562592331;
array[4593]=30'd919054939;
array[4594]=30'd898043496;
array[4595]=30'd919054939;
array[4596]=30'd898043496;
array[4597]=30'd898043496;
array[4598]=30'd919054939;
array[4599]=30'd898043496;
array[4600]=30'd919054939;
array[4601]=30'd898043496;
array[4602]=30'd919054939;
array[4603]=30'd919054939;
array[4604]=30'd919054939;
array[4605]=30'd919054939;
array[4606]=30'd919054939;
array[4607]=30'd919054939;
array[4608]=30'd898043496;
array[4609]=30'd919054939;
array[4610]=30'd919054939;
array[4611]=30'd919054939;
array[4612]=30'd919054939;
array[4613]=30'd919054939;
array[4614]=30'd919054939;
array[4615]=30'd919054939;
array[4616]=30'd919054939;
array[4617]=30'd919054939;
array[4618]=30'd919054939;
array[4619]=30'd919054939;
array[4620]=30'd919054939;
array[4621]=30'd919054939;
array[4622]=30'd919054939;
array[4623]=30'd919054939;
array[4624]=30'd842499661;
array[4625]=30'd795279924;
array[4626]=30'd979842606;
array[4627]=30'd959928886;
array[4628]=30'd959928886;
array[4629]=30'd979842606;
array[4630]=30'd979842606;
array[4631]=30'd959928886;
array[4632]=30'd959928886;
array[4633]=30'd959928886;
array[4634]=30'd795279924;
array[4635]=30'd938933826;
array[4636]=30'd919054939;
array[4637]=30'd919054939;
array[4638]=30'd919054939;
array[4639]=30'd919054939;
array[4640]=30'd919054939;
array[4641]=30'd919054939;
array[4642]=30'd919054939;
array[4643]=30'd919054939;
array[4644]=30'd919054939;
array[4645]=30'd919054939;
array[4646]=30'd884420162;
array[4647]=30'd482898518;
array[4648]=30'd478743092;
array[4649]=30'd473528913;
array[4650]=30'd473528913;
array[4651]=30'd461984322;
array[4652]=30'd391685709;
array[4653]=30'd300459585;
array[4654]=30'd421031501;
array[4655]=30'd473528913;
array[4656]=30'd473528913;
array[4657]=30'd488205898;
array[4658]=30'd488205898;
array[4659]=30'd488205898;
array[4660]=30'd488205898;
array[4661]=30'd473528913;
array[4662]=30'd473528913;
array[4663]=30'd461984322;
array[4664]=30'd434727495;
array[4665]=30'd488205898;
array[4666]=30'd488205898;
array[4667]=30'd488205898;
array[4668]=30'd488205898;
array[4669]=30'd488205898;
array[4670]=30'd473528913;
array[4671]=30'd488205898;
array[4672]=30'd461984322;
array[4673]=30'd373855782;
array[4674]=30'd300459585;
array[4675]=30'd452485730;
array[4676]=30'd461984322;
array[4677]=30'd461984322;
array[4678]=30'd314134080;
array[4679]=30'd461984322;
array[4680]=30'd461984322;
array[4681]=30'd370760263;
array[4682]=30'd473528913;
array[4683]=30'd461984322;
array[4684]=30'd473528913;
array[4685]=30'd473528913;
array[4686]=30'd473528913;
array[4687]=30'd461984322;
array[4688]=30'd482898518;
array[4689]=30'd898098744;
array[4690]=30'd919054939;
array[4691]=30'd919054939;
array[4692]=30'd919054939;
array[4693]=30'd919054939;
array[4694]=30'd919054939;
array[4695]=30'd919054939;
array[4696]=30'd919054939;
array[4697]=30'd919054939;
array[4698]=30'd959928886;
array[4699]=30'd936883742;
array[4700]=30'd877139478;
array[4701]=30'd877139478;
array[4702]=30'd898098744;
array[4703]=30'd959928886;
array[4704]=30'd919054939;
array[4705]=30'd919054939;
array[4706]=30'd919054939;
array[4707]=30'd919054939;
array[4708]=30'd919054939;
array[4709]=30'd919054939;
array[4710]=30'd919054939;
array[4711]=30'd919054939;
array[4712]=30'd919054939;
array[4713]=30'd919054939;
array[4714]=30'd919054939;
array[4715]=30'd919054939;
array[4716]=30'd919054939;
array[4717]=30'd919054939;
array[4718]=30'd919054939;
array[4719]=30'd919054939;
array[4720]=30'd919054939;
array[4721]=30'd725052963;
array[4722]=30'd959928886;
array[4723]=30'd959928886;
array[4724]=30'd959928886;
array[4725]=30'd959928886;
array[4726]=30'd979842606;
array[4727]=30'd959928886;
array[4728]=30'd959928886;
array[4729]=30'd959928886;
array[4730]=30'd694642226;
array[4731]=30'd938933826;
array[4732]=30'd938933826;
array[4733]=30'd919054939;
array[4734]=30'd919054939;
array[4735]=30'd919054939;
array[4736]=30'd919054939;
array[4737]=30'd919054939;
array[4738]=30'd919054939;
array[4739]=30'd919054939;
array[4740]=30'd919054939;
array[4741]=30'd919054939;
array[4742]=30'd562592331;
array[4743]=30'd482898518;
array[4744]=30'd473528913;
array[4745]=30'd488205898;
array[4746]=30'd488205898;
array[4747]=30'd488205898;
array[4748]=30'd370760263;
array[4749]=30'd335057455;
array[4750]=30'd391685709;
array[4751]=30'd473528913;
array[4752]=30'd473528913;
array[4753]=30'd488205898;
array[4754]=30'd488205898;
array[4755]=30'd488205898;
array[4756]=30'd488205898;
array[4757]=30'd473528913;
array[4758]=30'd473528913;
array[4759]=30'd370760263;
array[4760]=30'd461984322;
array[4761]=30'd473528913;
array[4762]=30'd488205898;
array[4763]=30'd488205898;
array[4764]=30'd473528913;
array[4765]=30'd488205898;
array[4766]=30'd488205898;
array[4767]=30'd473528913;
array[4768]=30'd461984322;
array[4769]=30'd370760263;
array[4770]=30'd252253768;
array[4771]=30'd461984322;
array[4772]=30'd473528913;
array[4773]=30'd473528913;
array[4774]=30'd461984322;
array[4775]=30'd434727495;
array[4776]=30'd434727495;
array[4777]=30'd434727495;
array[4778]=30'd473528913;
array[4779]=30'd473528913;
array[4780]=30'd473528913;
array[4781]=30'd473528913;
array[4782]=30'd473528913;
array[4783]=30'd473528913;
array[4784]=30'd421031501;
array[4785]=30'd842499661;
array[4786]=30'd919054939;
array[4787]=30'd919054939;
array[4788]=30'd919054939;
array[4789]=30'd919054939;
array[4790]=30'd919054939;
array[4791]=30'd959928886;
array[4792]=30'd936883742;
array[4793]=30'd857224695;
array[4794]=30'd833115609;
array[4795]=30'd798493124;
array[4796]=30'd774396326;
array[4797]=30'd758671804;
array[4798]=30'd785935846;
array[4799]=30'd898119130;
array[4800]=30'd877139478;
array[4801]=30'd936883742;
array[4802]=30'd919054939;
array[4803]=30'd919054939;
array[4804]=30'd919054939;
array[4805]=30'd919054939;
array[4806]=30'd919054939;
array[4807]=30'd919054939;
array[4808]=30'd919054939;
array[4809]=30'd919054939;
array[4810]=30'd919054939;
array[4811]=30'd919054939;
array[4812]=30'd919054939;
array[4813]=30'd919054939;
array[4814]=30'd919054939;
array[4815]=30'd919054939;
array[4816]=30'd919054939;
array[4817]=30'd779606588;
array[4818]=30'd916921900;
array[4819]=30'd959928886;
array[4820]=30'd979842606;
array[4821]=30'd959928886;
array[4822]=30'd959928886;
array[4823]=30'd959928886;
array[4824]=30'd959928886;
array[4825]=30'd959928886;
array[4826]=30'd555187752;
array[4827]=30'd884420162;
array[4828]=30'd919054939;
array[4829]=30'd919054939;
array[4830]=30'd919054939;
array[4831]=30'd919054939;
array[4832]=30'd919054939;
array[4833]=30'd919054939;
array[4834]=30'd919054939;
array[4835]=30'd919054939;
array[4836]=30'd919054939;
array[4837]=30'd656960070;
array[4838]=30'd482898518;
array[4839]=30'd473528913;
array[4840]=30'd473528913;
array[4841]=30'd488205898;
array[4842]=30'd488205898;
array[4843]=30'd461984322;
array[4844]=30'd434727495;
array[4845]=30'd461984322;
array[4846]=30'd346647116;
array[4847]=30'd461984322;
array[4848]=30'd473528913;
array[4849]=30'd473528913;
array[4850]=30'd488205898;
array[4851]=30'd473528913;
array[4852]=30'd473528913;
array[4853]=30'd473528913;
array[4854]=30'd461984322;
array[4855]=30'd370760263;
array[4856]=30'd473528913;
array[4857]=30'd473528913;
array[4858]=30'd473528913;
array[4859]=30'd473528913;
array[4860]=30'd473528913;
array[4861]=30'd488205898;
array[4862]=30'd473528913;
array[4863]=30'd473528913;
array[4864]=30'd461984322;
array[4865]=30'd482898518;
array[4866]=30'd335057455;
array[4867]=30'd478743092;
array[4868]=30'd461984322;
array[4869]=30'd473528913;
array[4870]=30'd473528913;
array[4871]=30'd461984322;
array[4872]=30'd370760263;
array[4873]=30'd473528913;
array[4874]=30'd473528913;
array[4875]=30'd473528913;
array[4876]=30'd473528913;
array[4877]=30'd473528913;
array[4878]=30'd473528913;
array[4879]=30'd473528913;
array[4880]=30'd434727495;
array[4881]=30'd725091917;
array[4882]=30'd919054939;
array[4883]=30'd919054939;
array[4884]=30'd919054939;
array[4885]=30'd919054939;
array[4886]=30'd959928886;
array[4887]=30'd983039487;
array[4888]=30'd785935846;
array[4889]=30'd758671804;
array[4890]=30'd774396326;
array[4891]=30'd790145435;
array[4892]=30'd885566856;
array[4893]=30'd850952611;
array[4894]=30'd774396326;
array[4895]=30'd816348600;
array[4896]=30'd833115609;
array[4897]=30'd921177592;
array[4898]=30'd936883742;
array[4899]=30'd877139478;
array[4900]=30'd898098744;
array[4901]=30'd919054939;
array[4902]=30'd919054939;
array[4903]=30'd919054939;
array[4904]=30'd919054939;
array[4905]=30'd919054939;
array[4906]=30'd919054939;
array[4907]=30'd919054939;
array[4908]=30'd919054939;
array[4909]=30'd919054939;
array[4910]=30'd919054939;
array[4911]=30'd919054939;
array[4912]=30'd919054939;
array[4913]=30'd898098744;
array[4914]=30'd756500033;
array[4915]=30'd979842606;
array[4916]=30'd979842606;
array[4917]=30'd959928886;
array[4918]=30'd959928886;
array[4919]=30'd979842606;
array[4920]=30'd959928886;
array[4921]=30'd916921900;
array[4922]=30'd694642226;
array[4923]=30'd756500033;
array[4924]=30'd959928886;
array[4925]=30'd919054939;
array[4926]=30'd919054939;
array[4927]=30'd919054939;
array[4928]=30'd919054939;
array[4929]=30'd919054939;
array[4930]=30'd919054939;
array[4931]=30'd919054939;
array[4932]=30'd656960070;
array[4933]=30'd482898518;
array[4934]=30'd488205898;
array[4935]=30'd473528913;
array[4936]=30'd488205898;
array[4937]=30'd488205898;
array[4938]=30'd461984322;
array[4939]=30'd434727495;
array[4940]=30'd473528913;
array[4941]=30'd473528913;
array[4942]=30'd473528913;
array[4943]=30'd461984322;
array[4944]=30'd473528913;
array[4945]=30'd473528913;
array[4946]=30'd473528913;
array[4947]=30'd473528913;
array[4948]=30'd473528913;
array[4949]=30'd461984322;
array[4950]=30'd370760263;
array[4951]=30'd461984322;
array[4952]=30'd473528913;
array[4953]=30'd473528913;
array[4954]=30'd473528913;
array[4955]=30'd473528913;
array[4956]=30'd488205898;
array[4957]=30'd473528913;
array[4958]=30'd473528913;
array[4959]=30'd473528913;
array[4960]=30'd542675507;
array[4961]=30'd810005031;
array[4962]=30'd641178190;
array[4963]=30'd656960070;
array[4964]=30'd478743092;
array[4965]=30'd461984322;
array[4966]=30'd473528913;
array[4967]=30'd461984322;
array[4968]=30'd314134080;
array[4969]=30'd434727495;
array[4970]=30'd434727495;
array[4971]=30'd461984322;
array[4972]=30'd473528913;
array[4973]=30'd473528913;
array[4974]=30'd473528913;
array[4975]=30'd473528913;
array[4976]=30'd461984322;
array[4977]=30'd542675507;
array[4978]=30'd919054939;
array[4979]=30'd919054939;
array[4980]=30'd919054939;
array[4981]=30'd959928886;
array[4982]=30'd1000848926;
array[4983]=30'd857224695;
array[4984]=30'd790145435;
array[4985]=30'd885566856;
array[4986]=30'd885566856;
array[4987]=30'd816348600;
array[4988]=30'd911766951;
array[4989]=30'd996684226;
array[4990]=30'd871910847;
array[4991]=30'd758671804;
array[4992]=30'd798493124;
array[4993]=30'd925360587;
array[4994]=30'd921177592;
array[4995]=30'd821544417;
array[4996]=30'd936883742;
array[4997]=30'd938933826;
array[4998]=30'd919054939;
array[4999]=30'd919054939;
array[5000]=30'd919054939;
array[5001]=30'd919054939;
array[5002]=30'd919054939;
array[5003]=30'd919054939;
array[5004]=30'd919054939;
array[5005]=30'd919054939;
array[5006]=30'd919054939;
array[5007]=30'd919054939;
array[5008]=30'd919054939;
array[5009]=30'd919054939;
array[5010]=30'd810005031;
array[5011]=30'd884420162;
array[5012]=30'd959928886;
array[5013]=30'd959928886;
array[5014]=30'd959928886;
array[5015]=30'd959928886;
array[5016]=30'd860309028;
array[5017]=30'd725052963;
array[5018]=30'd936883742;
array[5019]=30'd860309028;
array[5020]=30'd842499661;
array[5021]=30'd919054939;
array[5022]=30'd919054939;
array[5023]=30'd919054939;
array[5024]=30'd919054939;
array[5025]=30'd919054939;
array[5026]=30'd919054939;
array[5027]=30'd725091917;
array[5028]=30'd482898518;
array[5029]=30'd473528913;
array[5030]=30'd473528913;
array[5031]=30'd473528913;
array[5032]=30'd488205898;
array[5033]=30'd473528913;
array[5034]=30'd434727495;
array[5035]=30'd473528913;
array[5036]=30'd473528913;
array[5037]=30'd488205898;
array[5038]=30'd488205898;
array[5039]=30'd488205898;
array[5040]=30'd473528913;
array[5041]=30'd488205898;
array[5042]=30'd473528913;
array[5043]=30'd473528913;
array[5044]=30'd370760263;
array[5045]=30'd370760263;
array[5046]=30'd370760263;
array[5047]=30'd473528913;
array[5048]=30'd473528913;
array[5049]=30'd473528913;
array[5050]=30'd473528913;
array[5051]=30'd473528913;
array[5052]=30'd473528913;
array[5053]=30'd473528913;
array[5054]=30'd473528913;
array[5055]=30'd524875335;
array[5056]=30'd842499661;
array[5057]=30'd641178190;
array[5058]=30'd694642226;
array[5059]=30'd641178190;
array[5060]=30'd478743092;
array[5061]=30'd461984322;
array[5062]=30'd461984322;
array[5063]=30'd434727495;
array[5064]=30'd810005031;
array[5065]=30'd936883742;
array[5066]=30'd898098744;
array[5067]=30'd542675507;
array[5068]=30'd461984322;
array[5069]=30'd473528913;
array[5070]=30'd473528913;
array[5071]=30'd473528913;
array[5072]=30'd473528913;
array[5073]=30'd478743092;
array[5074]=30'd725091917;
array[5075]=30'd919054939;
array[5076]=30'd919054939;
array[5077]=30'd979842606;
array[5078]=30'd921177592;
array[5079]=30'd774396326;
array[5080]=30'd850952611;
array[5081]=30'd911766951;
array[5082]=30'd790145435;
array[5083]=30'd740853147;
array[5084]=30'd816348600;
array[5085]=30'd996684226;
array[5086]=30'd911766951;
array[5087]=30'd774396326;
array[5088]=30'd798493124;
array[5089]=30'd925360587;
array[5090]=30'd964180446;
array[5091]=30'd785935846;
array[5092]=30'd903304711;
array[5093]=30'd916921900;
array[5094]=30'd919054939;
array[5095]=30'd919054939;
array[5096]=30'd919054939;
array[5097]=30'd919054939;
array[5098]=30'd919054939;
array[5099]=30'd919054939;
array[5100]=30'd919054939;
array[5101]=30'd919054939;
array[5102]=30'd919054939;
array[5103]=30'd919054939;
array[5104]=30'd919054939;
array[5105]=30'd919054939;
array[5106]=30'd919054939;
array[5107]=30'd779606588;
array[5108]=30'd779606588;
array[5109]=30'd756500033;
array[5110]=30'd668430907;
array[5111]=30'd649571855;
array[5112]=30'd649571855;
array[5113]=30'd903304711;
array[5114]=30'd959928886;
array[5115]=30'd959928886;
array[5116]=30'd795279924;
array[5117]=30'd884420162;
array[5118]=30'd919054939;
array[5119]=30'd919054939;
array[5120]=30'd919054939;
array[5121]=30'd919054939;
array[5122]=30'd725091917;
array[5123]=30'd482898518;
array[5124]=30'd473528913;
array[5125]=30'd473528913;
array[5126]=30'd488205898;
array[5127]=30'd488205898;
array[5128]=30'd488205898;
array[5129]=30'd434727495;
array[5130]=30'd461984322;
array[5131]=30'd473528913;
array[5132]=30'd473528913;
array[5133]=30'd488205898;
array[5134]=30'd488205898;
array[5135]=30'd488205898;
array[5136]=30'd488205898;
array[5137]=30'd488205898;
array[5138]=30'd473528913;
array[5139]=30'd473528913;
array[5140]=30'd434727495;
array[5141]=30'd370760263;
array[5142]=30'd434727495;
array[5143]=30'd473528913;
array[5144]=30'd473528913;
array[5145]=30'd473528913;
array[5146]=30'd473528913;
array[5147]=30'd473528913;
array[5148]=30'd473528913;
array[5149]=30'd473528913;
array[5150]=30'd488205898;
array[5151]=30'd524875335;
array[5152]=30'd702044720;
array[5153]=30'd756500033;
array[5154]=30'd795279924;
array[5155]=30'd725052963;
array[5156]=30'd490215960;
array[5157]=30'd478743092;
array[5158]=30'd490215960;
array[5159]=30'd490215960;
array[5160]=30'd810005031;
array[5161]=30'd779606588;
array[5162]=30'd810005031;
array[5163]=30'd584602166;
array[5164]=30'd444087878;
array[5165]=30'd461984322;
array[5166]=30'd473528913;
array[5167]=30'd473528913;
array[5168]=30'd473528913;
array[5169]=30'd461984322;
array[5170]=30'd421031501;
array[5171]=30'd842499661;
array[5172]=30'd979842606;
array[5173]=30'd1000848926;
array[5174]=30'd833115609;
array[5175]=30'd774396326;
array[5176]=30'd885566856;
array[5177]=30'd763929993;
array[5178]=30'd790145435;
array[5179]=30'd832088453;
array[5180]=30'd790145435;
array[5181]=30'd945316283;
array[5182]=30'd911766951;
array[5183]=30'd758671804;
array[5184]=30'd852917899;
array[5185]=30'd852917899;
array[5186]=30'd852917899;
array[5187]=30'd852917899;
array[5188]=30'd852917899;
array[5189]=30'd852917899;
array[5190]=30'd852917899;
array[5191]=30'd852917899;
array[5192]=30'd852917899;
array[5193]=30'd852917899;
array[5194]=30'd852917899;
array[5195]=30'd852917899;
array[5196]=30'd852917899;
array[5197]=30'd852917899;
array[5198]=30'd852917899;
array[5199]=30'd852917899;
array[5200]=30'd852917899;
array[5201]=30'd852917899;
array[5202]=30'd852917899;
array[5203]=30'd852917899;
array[5204]=30'd852917899;
array[5205]=30'd852917899;
array[5206]=30'd852917899;
array[5207]=30'd852917899;
array[5208]=30'd852917899;
array[5209]=30'd852917899;
array[5210]=30'd873911932;
array[5211]=30'd900139626;
array[5212]=30'd898096696;
array[5213]=30'd855119352;
array[5214]=30'd832058842;
array[5215]=30'd832058842;
array[5216]=30'd842495488;
array[5217]=30'd884422147;
array[5218]=30'd820432476;
array[5219]=30'd820432476;
array[5220]=30'd852917899;
array[5221]=30'd852917899;
array[5222]=30'd852917899;
array[5223]=30'd852917899;
array[5224]=30'd852917899;
array[5225]=30'd852917899;
array[5226]=30'd852917899;
array[5227]=30'd734429821;
array[5228]=30'd461756049;
array[5229]=30'd496374434;
array[5230]=30'd553991871;
array[5231]=30'd608524977;
array[5232]=30'd608524977;
array[5233]=30'd525668044;
array[5234]=30'd644157123;
array[5235]=30'd644157123;
array[5236]=30'd581260986;
array[5237]=30'd581260986;
array[5238]=30'd629468885;
array[5239]=30'd629468885;
array[5240]=30'd608524977;
array[5241]=30'd650530435;
array[5242]=30'd525726362;
array[5243]=30'd661993129;
array[5244]=30'd629468885;
array[5245]=30'd629468885;
array[5246]=30'd629468885;
array[5247]=30'd629468885;
array[5248]=30'd629468885;
array[5249]=30'd629468885;
array[5250]=30'd644157123;
array[5251]=30'd629468885;
array[5252]=30'd629468885;
array[5253]=30'd581260986;
array[5254]=30'd362128040;
array[5255]=30'd608524977;
array[5256]=30'd644157123;
array[5257]=30'd629468885;
array[5258]=30'd629468885;
array[5259]=30'd629468885;
array[5260]=30'd629468885;
array[5261]=30'd629468885;
array[5262]=30'd644157123;
array[5263]=30'd615902883;
array[5264]=30'd815162003;
array[5265]=30'd852917899;
array[5266]=30'd815162003;
array[5267]=30'd815162003;
array[5268]=30'd815162003;
array[5269]=30'd852917899;
array[5270]=30'd815162003;
array[5271]=30'd852917899;
array[5272]=30'd852917899;
array[5273]=30'd852917899;
array[5274]=30'd852917899;
array[5275]=30'd852917899;
array[5276]=30'd852917899;
array[5277]=30'd852917899;
array[5278]=30'd852917899;
array[5279]=30'd873911932;
array[5280]=30'd852917899;
array[5281]=30'd852917899;
array[5282]=30'd852917899;
array[5283]=30'd852917899;
array[5284]=30'd852917899;
array[5285]=30'd852917899;
array[5286]=30'd852917899;
array[5287]=30'd852917899;
array[5288]=30'd852917899;
array[5289]=30'd852917899;
array[5290]=30'd852917899;
array[5291]=30'd852917899;
array[5292]=30'd852917899;
array[5293]=30'd852917899;
array[5294]=30'd852917899;
array[5295]=30'd852917899;
array[5296]=30'd852917899;
array[5297]=30'd852917899;
array[5298]=30'd852917899;
array[5299]=30'd852917899;
array[5300]=30'd852917899;
array[5301]=30'd852917899;
array[5302]=30'd852917899;
array[5303]=30'd852917899;
array[5304]=30'd852917899;
array[5305]=30'd852917899;
array[5306]=30'd852917899;
array[5307]=30'd873911932;
array[5308]=30'd884420162;
array[5309]=30'd916923947;
array[5310]=30'd884422147;
array[5311]=30'd884422147;
array[5312]=30'd860306981;
array[5313]=30'd884420162;
array[5314]=30'd873911932;
array[5315]=30'd852917899;
array[5316]=30'd852917899;
array[5317]=30'd852917899;
array[5318]=30'd852917899;
array[5319]=30'd852917899;
array[5320]=30'd852917899;
array[5321]=30'd852917899;
array[5322]=30'd815162003;
array[5323]=30'd559296136;
array[5324]=30'd496374434;
array[5325]=30'd591795877;
array[5326]=30'd444952244;
array[5327]=30'd608524977;
array[5328]=30'd516257448;
array[5329]=30'd608524977;
array[5330]=30'd644157123;
array[5331]=30'd644157123;
array[5332]=30'd485848753;
array[5333]=30'd644157123;
array[5334]=30'd629468885;
array[5335]=30'd644157123;
array[5336]=30'd548772504;
array[5337]=30'd820432476;
array[5338]=30'd530993763;
array[5339]=30'd661993129;
array[5340]=30'd629468885;
array[5341]=30'd629468885;
array[5342]=30'd629468885;
array[5343]=30'd629468885;
array[5344]=30'd629468885;
array[5345]=30'd629468885;
array[5346]=30'd644157123;
array[5347]=30'd629468885;
array[5348]=30'd629468885;
array[5349]=30'd644157123;
array[5350]=30'd394645149;
array[5351]=30'd496374434;
array[5352]=30'd661993129;
array[5353]=30'd644157123;
array[5354]=30'd629468885;
array[5355]=30'd629468885;
array[5356]=30'd644157123;
array[5357]=30'd629468885;
array[5358]=30'd644157123;
array[5359]=30'd581260986;
array[5360]=30'd650530435;
array[5361]=30'd791076458;
array[5362]=30'd820432476;
array[5363]=30'd852917899;
array[5364]=30'd852917899;
array[5365]=30'd852917899;
array[5366]=30'd852917899;
array[5367]=30'd815162003;
array[5368]=30'd852917899;
array[5369]=30'd852917899;
array[5370]=30'd852917899;
array[5371]=30'd852917899;
array[5372]=30'd852917899;
array[5373]=30'd852917899;
array[5374]=30'd873911932;
array[5375]=30'd900139626;
array[5376]=30'd852917899;
array[5377]=30'd852917899;
array[5378]=30'd852917899;
array[5379]=30'd852917899;
array[5380]=30'd852917899;
array[5381]=30'd852917899;
array[5382]=30'd852917899;
array[5383]=30'd852917899;
array[5384]=30'd852917899;
array[5385]=30'd852917899;
array[5386]=30'd852917899;
array[5387]=30'd852917899;
array[5388]=30'd852917899;
array[5389]=30'd852917899;
array[5390]=30'd852917899;
array[5391]=30'd852917899;
array[5392]=30'd852917899;
array[5393]=30'd852917899;
array[5394]=30'd852917899;
array[5395]=30'd852917899;
array[5396]=30'd852917899;
array[5397]=30'd852917899;
array[5398]=30'd852917899;
array[5399]=30'd852917899;
array[5400]=30'd852917899;
array[5401]=30'd852917899;
array[5402]=30'd852917899;
array[5403]=30'd852917899;
array[5404]=30'd873911932;
array[5405]=30'd873911932;
array[5406]=30'd884420162;
array[5407]=30'd839339599;
array[5408]=30'd839339599;
array[5409]=30'd852917899;
array[5410]=30'd852917899;
array[5411]=30'd852917899;
array[5412]=30'd852917899;
array[5413]=30'd852917899;
array[5414]=30'd852917899;
array[5415]=30'd852917899;
array[5416]=30'd852917899;
array[5417]=30'd852917899;
array[5418]=30'd777409151;
array[5419]=30'd496374434;
array[5420]=30'd461756049;
array[5421]=30'd634745492;
array[5422]=30'd485848753;
array[5423]=30'd661993129;
array[5424]=30'd485848753;
array[5425]=30'd661993129;
array[5426]=30'd644157123;
array[5427]=30'd608524977;
array[5428]=30'd516257448;
array[5429]=30'd644157123;
array[5430]=30'd629468885;
array[5431]=30'd591795877;
array[5432]=30'd791076458;
array[5433]=30'd839339599;
array[5434]=30'd530993763;
array[5435]=30'd661993129;
array[5436]=30'd629468885;
array[5437]=30'd629468885;
array[5438]=30'd629468885;
array[5439]=30'd629468885;
array[5440]=30'd644157123;
array[5441]=30'd629468885;
array[5442]=30'd644157123;
array[5443]=30'd629468885;
array[5444]=30'd629468885;
array[5445]=30'd629468885;
array[5446]=30'd516257448;
array[5447]=30'd368466587;
array[5448]=30'd661993129;
array[5449]=30'd629468885;
array[5450]=30'd629468885;
array[5451]=30'd629468885;
array[5452]=30'd525668044;
array[5453]=30'd608524977;
array[5454]=30'd644157123;
array[5455]=30'd661993129;
array[5456]=30'd559296136;
array[5457]=30'd852917899;
array[5458]=30'd820432476;
array[5459]=30'd852917899;
array[5460]=30'd815162003;
array[5461]=30'd815162003;
array[5462]=30'd852917899;
array[5463]=30'd852917899;
array[5464]=30'd852917899;
array[5465]=30'd852917899;
array[5466]=30'd852917899;
array[5467]=30'd852917899;
array[5468]=30'd873911932;
array[5469]=30'd900139626;
array[5470]=30'd941029952;
array[5471]=30'd963075636;
array[5472]=30'd852917899;
array[5473]=30'd852917899;
array[5474]=30'd852917899;
array[5475]=30'd852917899;
array[5476]=30'd852917899;
array[5477]=30'd852917899;
array[5478]=30'd852917899;
array[5479]=30'd852917899;
array[5480]=30'd852917899;
array[5481]=30'd852917899;
array[5482]=30'd852917899;
array[5483]=30'd852917899;
array[5484]=30'd852917899;
array[5485]=30'd852917899;
array[5486]=30'd852917899;
array[5487]=30'd852917899;
array[5488]=30'd852917899;
array[5489]=30'd852917899;
array[5490]=30'd852917899;
array[5491]=30'd852917899;
array[5492]=30'd852917899;
array[5493]=30'd852917899;
array[5494]=30'd852917899;
array[5495]=30'd852917899;
array[5496]=30'd852917899;
array[5497]=30'd852917899;
array[5498]=30'd852917899;
array[5499]=30'd852917899;
array[5500]=30'd852917899;
array[5501]=30'd852917899;
array[5502]=30'd852917899;
array[5503]=30'd852917899;
array[5504]=30'd852917899;
array[5505]=30'd852917899;
array[5506]=30'd852917899;
array[5507]=30'd852917899;
array[5508]=30'd852917899;
array[5509]=30'd852917899;
array[5510]=30'd852917899;
array[5511]=30'd852917899;
array[5512]=30'd852917899;
array[5513]=30'd852917899;
array[5514]=30'd650530435;
array[5515]=30'd496374434;
array[5516]=30'd591795877;
array[5517]=30'd553991871;
array[5518]=30'd553991871;
array[5519]=30'd608524977;
array[5520]=30'd516257448;
array[5521]=30'd644157123;
array[5522]=30'd644157123;
array[5523]=30'd516257448;
array[5524]=30'd548772504;
array[5525]=30'd629468885;
array[5526]=30'd644157123;
array[5527]=30'd582345342;
array[5528]=30'd941029952;
array[5529]=30'd839339599;
array[5530]=30'd556154453;
array[5531]=30'd634745492;
array[5532]=30'd581260986;
array[5533]=30'd644157123;
array[5534]=30'd629468885;
array[5535]=30'd608524977;
array[5536]=30'd525668044;
array[5537]=30'd629468885;
array[5538]=30'd629468885;
array[5539]=30'd629468885;
array[5540]=30'd629468885;
array[5541]=30'd629468885;
array[5542]=30'd553991871;
array[5543]=30'd300284569;
array[5544]=30'd591795877;
array[5545]=30'd629468885;
array[5546]=30'd629468885;
array[5547]=30'd629468885;
array[5548]=30'd629468885;
array[5549]=30'd525668044;
array[5550]=30'd644157123;
array[5551]=30'd644157123;
array[5552]=30'd548772504;
array[5553]=30'd777409151;
array[5554]=30'd852917899;
array[5555]=30'd852917899;
array[5556]=30'd852917899;
array[5557]=30'd852917899;
array[5558]=30'd852917899;
array[5559]=30'd852917899;
array[5560]=30'd852917899;
array[5561]=30'd852917899;
array[5562]=30'd852917899;
array[5563]=30'd873911932;
array[5564]=30'd920102487;
array[5565]=30'd963075636;
array[5566]=30'd915924476;
array[5567]=30'd832058842;
array[5568]=30'd852917899;
array[5569]=30'd852917899;
array[5570]=30'd852917899;
array[5571]=30'd852917899;
array[5572]=30'd852917899;
array[5573]=30'd852917899;
array[5574]=30'd852917899;
array[5575]=30'd852917899;
array[5576]=30'd852917899;
array[5577]=30'd852917899;
array[5578]=30'd852917899;
array[5579]=30'd852917899;
array[5580]=30'd852917899;
array[5581]=30'd852917899;
array[5582]=30'd852917899;
array[5583]=30'd852917899;
array[5584]=30'd852917899;
array[5585]=30'd852917899;
array[5586]=30'd852917899;
array[5587]=30'd873911932;
array[5588]=30'd873911932;
array[5589]=30'd852917899;
array[5590]=30'd852917899;
array[5591]=30'd852917899;
array[5592]=30'd852917899;
array[5593]=30'd852917899;
array[5594]=30'd852917899;
array[5595]=30'd852917899;
array[5596]=30'd852917899;
array[5597]=30'd852917899;
array[5598]=30'd852917899;
array[5599]=30'd852917899;
array[5600]=30'd852917899;
array[5601]=30'd852917899;
array[5602]=30'd852917899;
array[5603]=30'd852917899;
array[5604]=30'd852917899;
array[5605]=30'd852917899;
array[5606]=30'd852917899;
array[5607]=30'd852917899;
array[5608]=30'd852917899;
array[5609]=30'd815162003;
array[5610]=30'd496374434;
array[5611]=30'd461756049;
array[5612]=30'd634745492;
array[5613]=30'd485848753;
array[5614]=30'd608524977;
array[5615]=30'd548772504;
array[5616]=30'd553991871;
array[5617]=30'd644157123;
array[5618]=30'd661993129;
array[5619]=30'd496374434;
array[5620]=30'd591795877;
array[5621]=30'd644157123;
array[5622]=30'd608524977;
array[5623]=30'd739680847;
array[5624]=30'd941029952;
array[5625]=30'd884420162;
array[5626]=30'd530993763;
array[5627]=30'd634745492;
array[5628]=30'd444952244;
array[5629]=30'd608524977;
array[5630]=30'd644157123;
array[5631]=30'd644157123;
array[5632]=30'd427157133;
array[5633]=30'd644157123;
array[5634]=30'd629468885;
array[5635]=30'd629468885;
array[5636]=30'd629468885;
array[5637]=30'd608524977;
array[5638]=30'd608524977;
array[5639]=30'd328601227;
array[5640]=30'd525726362;
array[5641]=30'd644157123;
array[5642]=30'd629468885;
array[5643]=30'd629468885;
array[5644]=30'd629468885;
array[5645]=30'd525668044;
array[5646]=30'd644157123;
array[5647]=30'd644157123;
array[5648]=30'd608524977;
array[5649]=30'd702982791;
array[5650]=30'd852917899;
array[5651]=30'd852917899;
array[5652]=30'd852917899;
array[5653]=30'd852917899;
array[5654]=30'd852917899;
array[5655]=30'd852917899;
array[5656]=30'd852917899;
array[5657]=30'd852917899;
array[5658]=30'd852917899;
array[5659]=30'd873911932;
array[5660]=30'd884420162;
array[5661]=30'd819475993;
array[5662]=30'd776468978;
array[5663]=30'd794287561;
array[5664]=30'd852917899;
array[5665]=30'd852917899;
array[5666]=30'd852917899;
array[5667]=30'd852917899;
array[5668]=30'd852917899;
array[5669]=30'd852917899;
array[5670]=30'd852917899;
array[5671]=30'd852917899;
array[5672]=30'd852917899;
array[5673]=30'd852917899;
array[5674]=30'd873911932;
array[5675]=30'd873911932;
array[5676]=30'd900139626;
array[5677]=30'd900139626;
array[5678]=30'd900139626;
array[5679]=30'd884420162;
array[5680]=30'd884420162;
array[5681]=30'd839339599;
array[5682]=30'd839339599;
array[5683]=30'd884420162;
array[5684]=30'd941029952;
array[5685]=30'd884420162;
array[5686]=30'd839339599;
array[5687]=30'd884420162;
array[5688]=30'd873911932;
array[5689]=30'd852917899;
array[5690]=30'd852917899;
array[5691]=30'd852917899;
array[5692]=30'd852917899;
array[5693]=30'd852917899;
array[5694]=30'd852917899;
array[5695]=30'd852917899;
array[5696]=30'd852917899;
array[5697]=30'd852917899;
array[5698]=30'd852917899;
array[5699]=30'd852917899;
array[5700]=30'd852917899;
array[5701]=30'd852917899;
array[5702]=30'd852917899;
array[5703]=30'd852917899;
array[5704]=30'd852917899;
array[5705]=30'd734429821;
array[5706]=30'd503733877;
array[5707]=30'd461756049;
array[5708]=30'd661993129;
array[5709]=30'd444952244;
array[5710]=30'd661993129;
array[5711]=30'd516257448;
array[5712]=30'd608524977;
array[5713]=30'd661993129;
array[5714]=30'd591795877;
array[5715]=30'd582345342;
array[5716]=30'd591795877;
array[5717]=30'd661993129;
array[5718]=30'd548772504;
array[5719]=30'd884420162;
array[5720]=30'd941029952;
array[5721]=30'd884420162;
array[5722]=30'd512140869;
array[5723]=30'd625322602;
array[5724]=30'd650530435;
array[5725]=30'd559296136;
array[5726]=30'd661993129;
array[5727]=30'd661993129;
array[5728]=30'd496374434;
array[5729]=30'd548772504;
array[5730]=30'd661993129;
array[5731]=30'd629468885;
array[5732]=30'd629468885;
array[5733]=30'd485848753;
array[5734]=30'd608524977;
array[5735]=30'd328601227;
array[5736]=30'd461756049;
array[5737]=30'd661993129;
array[5738]=30'd629468885;
array[5739]=30'd629468885;
array[5740]=30'd629468885;
array[5741]=30'd608524977;
array[5742]=30'd553991871;
array[5743]=30'd644157123;
array[5744]=30'd661993129;
array[5745]=30'd591795877;
array[5746]=30'd852917899;
array[5747]=30'd852917899;
array[5748]=30'd852917899;
array[5749]=30'd852917899;
array[5750]=30'd852917899;
array[5751]=30'd852917899;
array[5752]=30'd852917899;
array[5753]=30'd852917899;
array[5754]=30'd852917899;
array[5755]=30'd852917899;
array[5756]=30'd873911932;
array[5757]=30'd839339599;
array[5758]=30'd808945195;
array[5759]=30'd842495488;
array[5760]=30'd852917899;
array[5761]=30'd852917899;
array[5762]=30'd852917899;
array[5763]=30'd852917899;
array[5764]=30'd852917899;
array[5765]=30'd852917899;
array[5766]=30'd852917899;
array[5767]=30'd852917899;
array[5768]=30'd852917899;
array[5769]=30'd873911932;
array[5770]=30'd900139626;
array[5771]=30'd920102487;
array[5772]=30'd936883742;
array[5773]=30'd875032088;
array[5774]=30'd819437027;
array[5775]=30'd794287561;
array[5776]=30'd794287561;
array[5777]=30'd794287561;
array[5778]=30'd776468978;
array[5779]=30'd842495488;
array[5780]=30'd963077644;
array[5781]=30'd855119352;
array[5782]=30'd808945195;
array[5783]=30'd860306981;
array[5784]=30'd839339599;
array[5785]=30'd852917899;
array[5786]=30'd852917899;
array[5787]=30'd852917899;
array[5788]=30'd852917899;
array[5789]=30'd852917899;
array[5790]=30'd852917899;
array[5791]=30'd852917899;
array[5792]=30'd852917899;
array[5793]=30'd852917899;
array[5794]=30'd852917899;
array[5795]=30'd852917899;
array[5796]=30'd852917899;
array[5797]=30'd852917899;
array[5798]=30'd852917899;
array[5799]=30'd852917899;
array[5800]=30'd820432476;
array[5801]=30'd559296136;
array[5802]=30'd559296136;
array[5803]=30'd496374434;
array[5804]=30'd661993129;
array[5805]=30'd485848753;
array[5806]=30'd661993129;
array[5807]=30'd461756049;
array[5808]=30'd608524977;
array[5809]=30'd661993129;
array[5810]=30'd559296136;
array[5811]=30'd739680847;
array[5812]=30'd604358258;
array[5813]=30'd661993129;
array[5814]=30'd650530435;
array[5815]=30'd941029952;
array[5816]=30'd941029952;
array[5817]=30'd941029952;
array[5818]=30'd512140869;
array[5819]=30'd604358258;
array[5820]=30'd756500033;
array[5821]=30'd530993763;
array[5822]=30'd634745492;
array[5823]=30'd661993129;
array[5824]=30'd650530435;
array[5825]=30'd589750888;
array[5826]=30'd634745492;
array[5827]=30'd644157123;
array[5828]=30'd644157123;
array[5829]=30'd444952244;
array[5830]=30'd591795877;
array[5831]=30'd374749802;
array[5832]=30'd368466587;
array[5833]=30'd661993129;
array[5834]=30'd629468885;
array[5835]=30'd629468885;
array[5836]=30'd629468885;
array[5837]=30'd644157123;
array[5838]=30'd516257448;
array[5839]=30'd644157123;
array[5840]=30'd644157123;
array[5841]=30'd548772504;
array[5842]=30'd852917899;
array[5843]=30'd852917899;
array[5844]=30'd852917899;
array[5845]=30'd852917899;
array[5846]=30'd852917899;
array[5847]=30'd852917899;
array[5848]=30'd852917899;
array[5849]=30'd852917899;
array[5850]=30'd852917899;
array[5851]=30'd852917899;
array[5852]=30'd852917899;
array[5853]=30'd873911932;
array[5854]=30'd873911932;
array[5855]=30'd884420162;
array[5856]=30'd852917899;
array[5857]=30'd852917899;
array[5858]=30'd852917899;
array[5859]=30'd852917899;
array[5860]=30'd852917899;
array[5861]=30'd852917899;
array[5862]=30'd852917899;
array[5863]=30'd852917899;
array[5864]=30'd873911932;
array[5865]=30'd873911932;
array[5866]=30'd941029952;
array[5867]=30'd963077644;
array[5868]=30'd832058842;
array[5869]=30'd764966339;
array[5870]=30'd834187654;
array[5871]=30'd790145435;
array[5872]=30'd810051001;
array[5873]=30'd810051001;
array[5874]=30'd764966339;
array[5875]=30'd794287561;
array[5876]=30'd884422147;
array[5877]=30'd915924476;
array[5878]=30'd776468978;
array[5879]=30'd819437027;
array[5880]=30'd860306981;
array[5881]=30'd873911932;
array[5882]=30'd852917899;
array[5883]=30'd852917899;
array[5884]=30'd852917899;
array[5885]=30'd852917899;
array[5886]=30'd852917899;
array[5887]=30'd852917899;
array[5888]=30'd852917899;
array[5889]=30'd852917899;
array[5890]=30'd852917899;
array[5891]=30'd852917899;
array[5892]=30'd852917899;
array[5893]=30'd852917899;
array[5894]=30'd852917899;
array[5895]=30'd852917899;
array[5896]=30'd839339599;
array[5897]=30'd484874837;
array[5898]=30'd559296136;
array[5899]=30'd548772504;
array[5900]=30'd661993129;
array[5901]=30'd452327079;
array[5902]=30'd608524977;
array[5903]=30'd368466587;
array[5904]=30'd634745492;
array[5905]=30'd608524977;
array[5906]=30'd589750888;
array[5907]=30'd793183798;
array[5908]=30'd582345342;
array[5909]=30'd634745492;
array[5910]=30'd739680847;
array[5911]=30'd963075636;
array[5912]=30'd941029952;
array[5913]=30'd941029952;
array[5914]=30'd664186439;
array[5915]=30'd589750888;
array[5916]=30'd820432476;
array[5917]=30'd756500033;
array[5918]=30'd582345342;
array[5919]=30'd661993129;
array[5920]=30'd568785526;
array[5921]=30'd756500033;
array[5922]=30'd582345342;
array[5923]=30'd661993129;
array[5924]=30'd644157123;
array[5925]=30'd548772504;
array[5926]=30'd525726362;
array[5927]=30'd433483392;
array[5928]=30'd374749802;
array[5929]=30'd634745492;
array[5930]=30'd644157123;
array[5931]=30'd629468885;
array[5932]=30'd629468885;
array[5933]=30'd629468885;
array[5934]=30'd516257448;
array[5935]=30'd644157123;
array[5936]=30'd644157123;
array[5937]=30'd548772504;
array[5938]=30'd815162003;
array[5939]=30'd852917899;
array[5940]=30'd852917899;
array[5941]=30'd852917899;
array[5942]=30'd852917899;
array[5943]=30'd852917899;
array[5944]=30'd852917899;
array[5945]=30'd852917899;
array[5946]=30'd852917899;
array[5947]=30'd852917899;
array[5948]=30'd852917899;
array[5949]=30'd852917899;
array[5950]=30'd852917899;
array[5951]=30'd900139626;
array[5952]=30'd852917899;
array[5953]=30'd852917899;
array[5954]=30'd852917899;
array[5955]=30'd852917899;
array[5956]=30'd852917899;
array[5957]=30'd852917899;
array[5958]=30'd873911932;
array[5959]=30'd873911932;
array[5960]=30'd873911932;
array[5961]=30'd920102487;
array[5962]=30'd1002945052;
array[5963]=30'd855119352;
array[5964]=30'd790145435;
array[5965]=30'd883468684;
array[5966]=30'd914919842;
array[5967]=30'd834187654;
array[5968]=30'd810051001;
array[5969]=30'd944268729;
array[5970]=30'd870853059;
array[5971]=30'd754446794;
array[5972]=30'd842495488;
array[5973]=30'd936883742;
array[5974]=30'd915924476;
array[5975]=30'd794287561;
array[5976]=30'd842495488;
array[5977]=30'd839339599;
array[5978]=30'd852917899;
array[5979]=30'd852917899;
array[5980]=30'd852917899;
array[5981]=30'd852917899;
array[5982]=30'd852917899;
array[5983]=30'd852917899;
array[5984]=30'd852917899;
array[5985]=30'd852917899;
array[5986]=30'd852917899;
array[5987]=30'd852917899;
array[5988]=30'd852917899;
array[5989]=30'd852917899;
array[5990]=30'd852917899;
array[5991]=30'd873911932;
array[5992]=30'd884420162;
array[5993]=30'd530993763;
array[5994]=30'd582345342;
array[5995]=30'd548772504;
array[5996]=30'd608524977;
array[5997]=30'd362128040;
array[5998]=30'd548772504;
array[5999]=30'd433483392;
array[6000]=30'd634745492;
array[6001]=30'd591795877;
array[6002]=30'd710361687;
array[6003]=30'd808945195;
array[6004]=30'd503733877;
array[6005]=30'd582345342;
array[6006]=30'd839339599;
array[6007]=30'd963075636;
array[6008]=30'd941029952;
array[6009]=30'd941029952;
array[6010]=30'd793183798;
array[6011]=30'd530993763;
array[6012]=30'd793183798;
array[6013]=30'd916923947;
array[6014]=30'd530993763;
array[6015]=30'd634745492;
array[6016]=30'd503733877;
array[6017]=30'd884420162;
array[6018]=30'd556154453;
array[6019]=30'd634745492;
array[6020]=30'd608524977;
array[6021]=30'd591795877;
array[6022]=30'd503733877;
array[6023]=30'd589750888;
array[6024]=30'd484874837;
array[6025]=30'd634745492;
array[6026]=30'd644157123;
array[6027]=30'd644157123;
array[6028]=30'd629468885;
array[6029]=30'd629468885;
array[6030]=30'd525668044;
array[6031]=30'd644157123;
array[6032]=30'd629468885;
array[6033]=30'd553991871;
array[6034]=30'd815162003;
array[6035]=30'd852917899;
array[6036]=30'd852917899;
array[6037]=30'd815162003;
array[6038]=30'd852917899;
array[6039]=30'd852917899;
array[6040]=30'd852917899;
array[6041]=30'd852917899;
array[6042]=30'd852917899;
array[6043]=30'd852917899;
array[6044]=30'd852917899;
array[6045]=30'd852917899;
array[6046]=30'd852917899;
array[6047]=30'd873911932;
array[6048]=30'd852917899;
array[6049]=30'd852917899;
array[6050]=30'd852917899;
array[6051]=30'd852917899;
array[6052]=30'd852917899;
array[6053]=30'd852917899;
array[6054]=30'd873911932;
array[6055]=30'd873911932;
array[6056]=30'd900139626;
array[6057]=30'd963075636;
array[6058]=30'd896012764;
array[6059]=30'd778588583;
array[6060]=30'd854099361;
array[6061]=30'd834187654;
array[6062]=30'd763929993;
array[6063]=30'd778588583;
array[6064]=30'd778588583;
array[6065]=30'd944268729;
array[6066]=30'd894973365;
array[6067]=30'd754446794;
array[6068]=30'd842495488;
array[6069]=30'd936883742;
array[6070]=30'd983039487;
array[6071]=30'd794287561;
array[6072]=30'd819437027;
array[6073]=30'd839339599;
array[6074]=30'd852917899;
array[6075]=30'd852917899;
array[6076]=30'd852917899;
array[6077]=30'd852917899;
array[6078]=30'd852917899;
array[6079]=30'd852917899;
array[6080]=30'd852917899;
array[6081]=30'd852917899;
array[6082]=30'd852917899;
array[6083]=30'd852917899;
array[6084]=30'd852917899;
array[6085]=30'd852917899;
array[6086]=30'd852917899;
array[6087]=30'd873911932;
array[6088]=30'd756500033;
array[6089]=30'd559296136;
array[6090]=30'd591795877;
array[6091]=30'd525726362;
array[6092]=30'd591795877;
array[6093]=30'd328601227;
array[6094]=30'd503733877;
array[6095]=30'd664186439;
array[6096]=30'd582345342;
array[6097]=30'd530993763;
array[6098]=30'd664186439;
array[6099]=30'd808945195;
array[6100]=30'd512140869;
array[6101]=30'd503733877;
array[6102]=30'd793183798;
array[6103]=30'd963075636;
array[6104]=30'd963075636;
array[6105]=30'd963075636;
array[6106]=30'd916923947;
array[6107]=30'd484874837;
array[6108]=30'd641178184;
array[6109]=30'd681011766;
array[6110]=30'd712433198;
array[6111]=30'd559296136;
array[6112]=30'd503733877;
array[6113]=30'd664186439;
array[6114]=30'd625394265;
array[6115]=30'd582345342;
array[6116]=30'd634745492;
array[6117]=30'd589750888;
array[6118]=30'd589750888;
array[6119]=30'd574048834;
array[6120]=30'd664186439;
array[6121]=30'd634745492;
array[6122]=30'd644157123;
array[6123]=30'd581260986;
array[6124]=30'd644157123;
array[6125]=30'd629468885;
array[6126]=30'd553991871;
array[6127]=30'd581260986;
array[6128]=30'd629468885;
array[6129]=30'd553991871;
array[6130]=30'd777409151;
array[6131]=30'd852917899;
array[6132]=30'd852917899;
array[6133]=30'd852917899;
array[6134]=30'd852917899;
array[6135]=30'd852917899;
array[6136]=30'd852917899;
array[6137]=30'd852917899;
array[6138]=30'd852917899;
array[6139]=30'd852917899;
array[6140]=30'd852917899;
array[6141]=30'd852917899;
array[6142]=30'd852917899;
array[6143]=30'd873911932;
array[6144]=30'd852917899;
array[6145]=30'd852917899;
array[6146]=30'd852917899;
array[6147]=30'd852917899;
array[6148]=30'd852917899;
array[6149]=30'd852917899;
array[6150]=30'd873911932;
array[6151]=30'd873911932;
array[6152]=30'd920102487;
array[6153]=30'd936883742;
array[6154]=30'd764966339;
array[6155]=30'd834187654;
array[6156]=30'd790145435;
array[6157]=30'd750292390;
array[6158]=30'd810051001;
array[6159]=30'd870853059;
array[6160]=30'd810051001;
array[6161]=30'd944268729;
array[6162]=30'd894973365;
array[6163]=30'd754446794;
array[6164]=30'd832058842;
array[6165]=30'd963077644;
array[6166]=30'd963129822;
array[6167]=30'd764966339;
array[6168]=30'd819437027;
array[6169]=30'd839339599;
array[6170]=30'd852917899;
array[6171]=30'd852917899;
array[6172]=30'd852917899;
array[6173]=30'd852917899;
array[6174]=30'd852917899;
array[6175]=30'd852917899;
array[6176]=30'd852917899;
array[6177]=30'd852917899;
array[6178]=30'd852917899;
array[6179]=30'd852917899;
array[6180]=30'd852917899;
array[6181]=30'd852917899;
array[6182]=30'd852917899;
array[6183]=30'd873911932;
array[6184]=30'd683036269;
array[6185]=30'd604358258;
array[6186]=30'd608524977;
array[6187]=30'd485848753;
array[6188]=30'd591795877;
array[6189]=30'd474371718;
array[6190]=30'd484874837;
array[6191]=30'd793183798;
array[6192]=30'd484874837;
array[6193]=30'd556154453;
array[6194]=30'd941029952;
array[6195]=30'd963075636;
array[6196]=30'd712433198;
array[6197]=30'd512140869;
array[6198]=30'd941029952;
array[6199]=30'd963075636;
array[6200]=30'd963075636;
array[6201]=30'd963075636;
array[6202]=30'd941029952;
array[6203]=30'd756500033;
array[6204]=30'd681011766;
array[6205]=30'd963075636;
array[6206]=30'd941029952;
array[6207]=30'd664186439;
array[6208]=30'd530993763;
array[6209]=30'd916923947;
array[6210]=30'd860306981;
array[6211]=30'd530993763;
array[6212]=30'd625322602;
array[6213]=30'd681011766;
array[6214]=30'd664186439;
array[6215]=30'd681011766;
array[6216]=30'd793183798;
array[6217]=30'd582345342;
array[6218]=30'd608524977;
array[6219]=30'd581260986;
array[6220]=30'd608524977;
array[6221]=30'd644157123;
array[6222]=30'd581260986;
array[6223]=30'd553991871;
array[6224]=30'd629468885;
array[6225]=30'd608524977;
array[6226]=30'd734429821;
array[6227]=30'd852917899;
array[6228]=30'd852917899;
array[6229]=30'd852917899;
array[6230]=30'd852917899;
array[6231]=30'd852917899;
array[6232]=30'd852917899;
array[6233]=30'd852917899;
array[6234]=30'd852917899;
array[6235]=30'd852917899;
array[6236]=30'd852917899;
array[6237]=30'd852917899;
array[6238]=30'd852917899;
array[6239]=30'd852917899;
array[6240]=30'd852917899;
array[6241]=30'd852917899;
array[6242]=30'd852917899;
array[6243]=30'd852917899;
array[6244]=30'd852917899;
array[6245]=30'd852917899;
array[6246]=30'd873911932;
array[6247]=30'd873911932;
array[6248]=30'd920102487;
array[6249]=30'd936883742;
array[6250]=30'd764966339;
array[6251]=30'd883468684;
array[6252]=30'd790145435;
array[6253]=30'd778588583;
array[6254]=30'd894973365;
array[6255]=30'd944268729;
array[6256]=30'd914919842;
array[6257]=30'd870853059;
array[6258]=30'd764966339;
array[6259]=30'd794287561;
array[6260]=30'd915924476;
array[6261]=30'd1002945052;
array[6262]=30'd855119352;
array[6263]=30'd794287561;
array[6264]=30'd842495488;
array[6265]=30'd839339599;
array[6266]=30'd852917899;
array[6267]=30'd852917899;
array[6268]=30'd852917899;
array[6269]=30'd852917899;
array[6270]=30'd852917899;
array[6271]=30'd852917899;
array[6272]=30'd852917899;
array[6273]=30'd852917899;
array[6274]=30'd852917899;
array[6275]=30'd852917899;
array[6276]=30'd852917899;
array[6277]=30'd852917899;
array[6278]=30'd873911932;
array[6279]=30'd873911932;
array[6280]=30'd625394265;
array[6281]=30'd634745492;
array[6282]=30'd661993129;
array[6283]=30'd444952244;
array[6284]=30'd548772504;
array[6285]=30'd674710128;
array[6286]=30'd421987917;
array[6287]=30'd712433198;
array[6288]=30'd580283972;
array[6289]=30'd547846737;
array[6290]=30'd963075636;
array[6291]=30'd963075636;
array[6292]=30'd884420162;
array[6293]=30'd574048834;
array[6294]=30'd963075636;
array[6295]=30'd963075636;
array[6296]=30'd963075636;
array[6297]=30'd963075636;
array[6298]=30'd963075636;
array[6299]=30'd941029952;
array[6300]=30'd793183798;
array[6301]=30'd981941808;
array[6302]=30'd963075636;
array[6303]=30'd884420162;
array[6304]=30'd528975414;
array[6305]=30'd916923947;
array[6306]=30'd963075636;
array[6307]=30'd739680847;
array[6308]=30'd484874837;
array[6309]=30'd756500033;
array[6310]=30'd724009508;
array[6311]=30'd756500033;
array[6312]=30'd756500033;
array[6313]=30'd484874837;
array[6314]=30'd634745492;
array[6315]=30'd553991871;
array[6316]=30'd608524977;
array[6317]=30'd644157123;
array[6318]=30'd608524977;
array[6319]=30'd525668044;
array[6320]=30'd629468885;
array[6321]=30'd608524977;
array[6322]=30'd702982791;
array[6323]=30'd852917899;
array[6324]=30'd852917899;
array[6325]=30'd852917899;
array[6326]=30'd852917899;
array[6327]=30'd852917899;
array[6328]=30'd852917899;
array[6329]=30'd852917899;
array[6330]=30'd852917899;
array[6331]=30'd852917899;
array[6332]=30'd852917899;
array[6333]=30'd852917899;
array[6334]=30'd852917899;
array[6335]=30'd852917899;
array[6336]=30'd852917899;
array[6337]=30'd852917899;
array[6338]=30'd852917899;
array[6339]=30'd852917899;
array[6340]=30'd852917899;
array[6341]=30'd873911932;
array[6342]=30'd873911932;
array[6343]=30'd873911932;
array[6344]=30'd900139626;
array[6345]=30'd936883742;
array[6346]=30'd764966339;
array[6347]=30'd810051001;
array[6348]=30'd894973365;
array[6349]=30'd778588583;
array[6350]=30'd810051001;
array[6351]=30'd894973365;
array[6352]=30'd810051001;
array[6353]=30'd764966339;
array[6354]=30'd810051001;
array[6355]=30'd896012764;
array[6356]=30'd963077644;
array[6357]=30'd963129822;
array[6358]=30'd764966339;
array[6359]=30'd819437027;
array[6360]=30'd860306981;
array[6361]=30'd873911932;
array[6362]=30'd852917899;
array[6363]=30'd852917899;
array[6364]=30'd852917899;
array[6365]=30'd852917899;
array[6366]=30'd852917899;
array[6367]=30'd852917899;
array[6368]=30'd852917899;
array[6369]=30'd852917899;
array[6370]=30'd852917899;
array[6371]=30'd852917899;
array[6372]=30'd852917899;
array[6373]=30'd852917899;
array[6374]=30'd873911932;
array[6375]=30'd852917899;
array[6376]=30'd589750888;
array[6377]=30'd634745492;
array[6378]=30'd661993129;
array[6379]=30'd516257448;
array[6380]=30'd525726362;
array[6381]=30'd739680847;
array[6382]=30'd470243883;
array[6383]=30'd916923947;
array[6384]=30'd860306981;
array[6385]=30'd574048834;
array[6386]=30'd963075636;
array[6387]=30'd963075636;
array[6388]=30'd963075636;
array[6389]=30'd916923947;
array[6390]=30'd963075636;
array[6391]=30'd963075636;
array[6392]=30'd963075636;
array[6393]=30'd963075636;
array[6394]=30'd963075636;
array[6395]=30'd963075636;
array[6396]=30'd963075636;
array[6397]=30'd963075636;
array[6398]=30'd963075636;
array[6399]=30'd963075636;
array[6400]=30'd884420162;
array[6401]=30'd941029952;
array[6402]=30'd963075636;
array[6403]=30'd884420162;
array[6404]=30'd512140869;
array[6405]=30'd839339599;
array[6406]=30'd598167087;
array[6407]=30'd808945195;
array[6408]=30'd445096449;
array[6409]=30'd503787028;
array[6410]=30'd456562280;
array[6411]=30'd525726362;
array[6412]=30'd608524977;
array[6413]=30'd644157123;
array[6414]=30'd644157123;
array[6415]=30'd553991871;
array[6416]=30'd644157123;
array[6417]=30'd581260986;
array[6418]=30'd734429821;
array[6419]=30'd852917899;
array[6420]=30'd852917899;
array[6421]=30'd852917899;
array[6422]=30'd852917899;
array[6423]=30'd852917899;
array[6424]=30'd852917899;
array[6425]=30'd852917899;
array[6426]=30'd852917899;
array[6427]=30'd852917899;
array[6428]=30'd852917899;
array[6429]=30'd852917899;
array[6430]=30'd852917899;
array[6431]=30'd852917899;
array[6432]=30'd852917899;
array[6433]=30'd852917899;
array[6434]=30'd852917899;
array[6435]=30'd852917899;
array[6436]=30'd852917899;
array[6437]=30'd852917899;
array[6438]=30'd873911932;
array[6439]=30'd873911932;
array[6440]=30'd900139626;
array[6441]=30'd936883742;
array[6442]=30'd855119352;
array[6443]=30'd764966339;
array[6444]=30'd896012764;
array[6445]=30'd870853059;
array[6446]=30'd764966339;
array[6447]=30'd764966339;
array[6448]=30'd794287561;
array[6449]=30'd842495488;
array[6450]=30'd875032088;
array[6451]=30'd936883742;
array[6452]=30'd983039487;
array[6453]=30'd832058842;
array[6454]=30'd819437027;
array[6455]=30'd860306981;
array[6456]=30'd839339599;
array[6457]=30'd852917899;
array[6458]=30'd852917899;
array[6459]=30'd852917899;
array[6460]=30'd852917899;
array[6461]=30'd852917899;
array[6462]=30'd852917899;
array[6463]=30'd852917899;
array[6464]=30'd852917899;
array[6465]=30'd852917899;
array[6466]=30'd852917899;
array[6467]=30'd852917899;
array[6468]=30'd873911932;
array[6469]=30'd873911932;
array[6470]=30'd852917899;
array[6471]=30'd852917899;
array[6472]=30'd568785526;
array[6473]=30'd661993129;
array[6474]=30'd661993129;
array[6475]=30'd608524977;
array[6476]=30'd427157133;
array[6477]=30'd756500033;
array[6478]=30'd860306981;
array[6479]=30'd963075636;
array[6480]=30'd963075636;
array[6481]=30'd884420162;
array[6482]=30'd963075636;
array[6483]=30'd963075636;
array[6484]=30'd963075636;
array[6485]=30'd963075636;
array[6486]=30'd963075636;
array[6487]=30'd963075636;
array[6488]=30'd963075636;
array[6489]=30'd963075636;
array[6490]=30'd963075636;
array[6491]=30'd963075636;
array[6492]=30'd963075636;
array[6493]=30'd963075636;
array[6494]=30'd963075636;
array[6495]=30'd963075636;
array[6496]=30'd963075636;
array[6497]=30'd963075636;
array[6498]=30'd963075636;
array[6499]=30'd963075636;
array[6500]=30'd916923947;
array[6501]=30'd963075636;
array[6502]=30'd860306981;
array[6503]=30'd808945195;
array[6504]=30'd650619404;
array[6505]=30'd819437027;
array[6506]=30'd450262593;
array[6507]=30'd503733877;
array[6508]=30'd634745492;
array[6509]=30'd644157123;
array[6510]=30'd644157123;
array[6511]=30'd553991871;
array[6512]=30'd644157123;
array[6513]=30'd581260986;
array[6514]=30'd777409151;
array[6515]=30'd852917899;
array[6516]=30'd852917899;
array[6517]=30'd852917899;
array[6518]=30'd852917899;
array[6519]=30'd852917899;
array[6520]=30'd852917899;
array[6521]=30'd852917899;
array[6522]=30'd852917899;
array[6523]=30'd852917899;
array[6524]=30'd852917899;
array[6525]=30'd852917899;
array[6526]=30'd852917899;
array[6527]=30'd852917899;
array[6528]=30'd852917899;
array[6529]=30'd852917899;
array[6530]=30'd852917899;
array[6531]=30'd852917899;
array[6532]=30'd852917899;
array[6533]=30'd873911932;
array[6534]=30'd873911932;
array[6535]=30'd873911932;
array[6536]=30'd873911932;
array[6537]=30'd900139626;
array[6538]=30'd936883742;
array[6539]=30'd776468978;
array[6540]=30'd794287561;
array[6541]=30'd855119352;
array[6542]=30'd832058842;
array[6543]=30'd819437027;
array[6544]=30'd884422147;
array[6545]=30'd898096696;
array[6546]=30'd936883742;
array[6547]=30'd983039487;
array[6548]=30'd896012764;
array[6549]=30'd794287561;
array[6550]=30'd842495488;
array[6551]=30'd839339599;
array[6552]=30'd852917899;
array[6553]=30'd852917899;
array[6554]=30'd852917899;
array[6555]=30'd852917899;
array[6556]=30'd852917899;
array[6557]=30'd852917899;
array[6558]=30'd852917899;
array[6559]=30'd852917899;
array[6560]=30'd852917899;
array[6561]=30'd852917899;
array[6562]=30'd852917899;
array[6563]=30'd852917899;
array[6564]=30'd852917899;
array[6565]=30'd852917899;
array[6566]=30'd873911932;
array[6567]=30'd852917899;
array[6568]=30'd559296136;
array[6569]=30'd634745492;
array[6570]=30'd608524977;
array[6571]=30'd581260986;
array[6572]=30'd525726362;
array[6573]=30'd756500033;
array[6574]=30'd963075636;
array[6575]=30'd963075636;
array[6576]=30'd963075636;
array[6577]=30'd963075636;
array[6578]=30'd884420162;
array[6579]=30'd884420162;
array[6580]=30'd916923947;
array[6581]=30'd963075636;
array[6582]=30'd963075636;
array[6583]=30'd963075636;
array[6584]=30'd963075636;
array[6585]=30'd963075636;
array[6586]=30'd963075636;
array[6587]=30'd963075636;
array[6588]=30'd963075636;
array[6589]=30'd963075636;
array[6590]=30'd963075636;
array[6591]=30'd963075636;
array[6592]=30'd963075636;
array[6593]=30'd963075636;
array[6594]=30'd963075636;
array[6595]=30'd963075636;
array[6596]=30'd963075636;
array[6597]=30'd963075636;
array[6598]=30'd963075636;
array[6599]=30'd875032088;
array[6600]=30'd650619404;
array[6601]=30'd776468978;
array[6602]=30'd512140869;
array[6603]=30'd484819572;
array[6604]=30'd634745492;
array[6605]=30'd644157123;
array[6606]=30'd644157123;
array[6607]=30'd553991871;
array[6608]=30'd644157123;
array[6609]=30'd553991871;
array[6610]=30'd777409151;
array[6611]=30'd852917899;
array[6612]=30'd852917899;
array[6613]=30'd852917899;
array[6614]=30'd852917899;
array[6615]=30'd852917899;
array[6616]=30'd852917899;
array[6617]=30'd852917899;
array[6618]=30'd852917899;
array[6619]=30'd852917899;
array[6620]=30'd852917899;
array[6621]=30'd852917899;
array[6622]=30'd852917899;
array[6623]=30'd852917899;
array[6624]=30'd852917899;
array[6625]=30'd852917899;
array[6626]=30'd852917899;
array[6627]=30'd852917899;
array[6628]=30'd852917899;
array[6629]=30'd873911932;
array[6630]=30'd873911932;
array[6631]=30'd873911932;
array[6632]=30'd873911932;
array[6633]=30'd900139626;
array[6634]=30'd920102487;
array[6635]=30'd855119352;
array[6636]=30'd764966339;
array[6637]=30'd832058842;
array[6638]=30'd896012764;
array[6639]=30'd915924476;
array[6640]=30'd915924476;
array[6641]=30'd915924476;
array[6642]=30'd896012764;
array[6643]=30'd832058842;
array[6644]=30'd785935846;
array[6645]=30'd819437027;
array[6646]=30'd860306981;
array[6647]=30'd873911932;
array[6648]=30'd852917899;
array[6649]=30'd852917899;
array[6650]=30'd852917899;
array[6651]=30'd852917899;
array[6652]=30'd852917899;
array[6653]=30'd852917899;
array[6654]=30'd852917899;
array[6655]=30'd852917899;
array[6656]=30'd852917899;
array[6657]=30'd852917899;
array[6658]=30'd852917899;
array[6659]=30'd852917899;
array[6660]=30'd852917899;
array[6661]=30'd852917899;
array[6662]=30'd852917899;
array[6663]=30'd852917899;
array[6664]=30'd582345342;
array[6665]=30'd634745492;
array[6666]=30'd661993129;
array[6667]=30'd485848753;
array[6668]=30'd615902883;
array[6669]=30'd756500033;
array[6670]=30'd963075636;
array[6671]=30'd963075636;
array[6672]=30'd860306981;
array[6673]=30'd724009508;
array[6674]=30'd724009508;
array[6675]=30'd860306981;
array[6676]=30'd808945195;
array[6677]=30'd808945195;
array[6678]=30'd963075636;
array[6679]=30'd981941808;
array[6680]=30'd963075636;
array[6681]=30'd963075636;
array[6682]=30'd963075636;
array[6683]=30'd963075636;
array[6684]=30'd963075636;
array[6685]=30'd916923947;
array[6686]=30'd808945195;
array[6687]=30'd724009508;
array[6688]=30'd724009508;
array[6689]=30'd756500033;
array[6690]=30'd916923947;
array[6691]=30'd963075636;
array[6692]=30'd963075636;
array[6693]=30'd963075636;
array[6694]=30'd963075636;
array[6695]=30'd860306981;
array[6696]=30'd503787028;
array[6697]=30'd470243883;
array[6698]=30'd556154453;
array[6699]=30'd484819572;
array[6700]=30'd608524977;
array[6701]=30'd644157123;
array[6702]=30'd608524977;
array[6703]=30'd553991871;
array[6704]=30'd629468885;
array[6705]=30'd516257448;
array[6706]=30'd815162003;
array[6707]=30'd852917899;
array[6708]=30'd852917899;
array[6709]=30'd852917899;
array[6710]=30'd852917899;
array[6711]=30'd852917899;
array[6712]=30'd852917899;
array[6713]=30'd852917899;
array[6714]=30'd852917899;
array[6715]=30'd852917899;
array[6716]=30'd852917899;
array[6717]=30'd852917899;
array[6718]=30'd852917899;
array[6719]=30'd852917899;
array[6720]=30'd852917899;
array[6721]=30'd873911932;
array[6722]=30'd873911932;
array[6723]=30'd852917899;
array[6724]=30'd873911932;
array[6725]=30'd873911932;
array[6726]=30'd873911932;
array[6727]=30'd873911932;
array[6728]=30'd873911932;
array[6729]=30'd873911932;
array[6730]=30'd884420162;
array[6731]=30'd898096696;
array[6732]=30'd855119352;
array[6733]=30'd764966339;
array[6734]=30'd778588583;
array[6735]=30'd764966339;
array[6736]=30'd778588583;
array[6737]=30'd778588583;
array[6738]=30'd778588583;
array[6739]=30'd794287561;
array[6740]=30'd842495488;
array[6741]=30'd860306981;
array[6742]=30'd839339599;
array[6743]=30'd873911932;
array[6744]=30'd852917899;
array[6745]=30'd852917899;
array[6746]=30'd852917899;
array[6747]=30'd852917899;
array[6748]=30'd852917899;
array[6749]=30'd873911932;
array[6750]=30'd873911932;
array[6751]=30'd852917899;
array[6752]=30'd873911932;
array[6753]=30'd873911932;
array[6754]=30'd873911932;
array[6755]=30'd873911932;
array[6756]=30'd873911932;
array[6757]=30'd873911932;
array[6758]=30'd852917899;
array[6759]=30'd852917899;
array[6760]=30'd589750888;
array[6761]=30'd634745492;
array[6762]=30'd661993129;
array[6763]=30'd485848753;
array[6764]=30'd666226344;
array[6765]=30'd625394265;
array[6766]=30'd898096696;
array[6767]=30'd756500033;
array[6768]=30'd756500033;
array[6769]=30'd756500033;
array[6770]=30'd470243883;
array[6771]=30'd336049694;
array[6772]=30'd598167087;
array[6773]=30'd916923947;
array[6774]=30'd963075636;
array[6775]=30'd963075636;
array[6776]=30'd981941808;
array[6777]=30'd963075636;
array[6778]=30'd963075636;
array[6779]=30'd963075636;
array[6780]=30'd941029952;
array[6781]=30'd756500033;
array[6782]=30'd808945195;
array[6783]=30'd724009508;
array[6784]=30'd681011766;
array[6785]=30'd724009508;
array[6786]=30'd681011766;
array[6787]=30'd724009508;
array[6788]=30'd916923947;
array[6789]=30'd963075636;
array[6790]=30'd963075636;
array[6791]=30'd936883742;
array[6792]=30'd724009508;
array[6793]=30'd530993763;
array[6794]=30'd625322602;
array[6795]=30'd452327079;
array[6796]=30'd644157123;
array[6797]=30'd644157123;
array[6798]=30'd608524977;
array[6799]=30'd525668044;
array[6800]=30'd644157123;
array[6801]=30'd548772504;
array[6802]=30'd852917899;
array[6803]=30'd852917899;
array[6804]=30'd852917899;
array[6805]=30'd852917899;
array[6806]=30'd852917899;
array[6807]=30'd852917899;
array[6808]=30'd852917899;
array[6809]=30'd852917899;
array[6810]=30'd852917899;
array[6811]=30'd852917899;
array[6812]=30'd852917899;
array[6813]=30'd852917899;
array[6814]=30'd852917899;
array[6815]=30'd852917899;
array[6816]=30'd852917899;
array[6817]=30'd873911932;
array[6818]=30'd873911932;
array[6819]=30'd873911932;
array[6820]=30'd873911932;
array[6821]=30'd873911932;
array[6822]=30'd873911932;
array[6823]=30'd873911932;
array[6824]=30'd873911932;
array[6825]=30'd873911932;
array[6826]=30'd900139626;
array[6827]=30'd898096696;
array[6828]=30'd915924476;
array[6829]=30'd832058842;
array[6830]=30'd819437027;
array[6831]=30'd819437027;
array[6832]=30'd819437027;
array[6833]=30'd842495488;
array[6834]=30'd842495488;
array[6835]=30'd860306981;
array[6836]=30'd860306981;
array[6837]=30'd884420162;
array[6838]=30'd873911932;
array[6839]=30'd873911932;
array[6840]=30'd852917899;
array[6841]=30'd852917899;
array[6842]=30'd873911932;
array[6843]=30'd873911932;
array[6844]=30'd873911932;
array[6845]=30'd873911932;
array[6846]=30'd873911932;
array[6847]=30'd873911932;
array[6848]=30'd873911932;
array[6849]=30'd873911932;
array[6850]=30'd873911932;
array[6851]=30'd873911932;
array[6852]=30'd873911932;
array[6853]=30'd852917899;
array[6854]=30'd852917899;
array[6855]=30'd873911932;
array[6856]=30'd625394265;
array[6857]=30'd634745492;
array[6858]=30'd661993129;
array[6859]=30'd485848753;
array[6860]=30'd666226344;
array[6861]=30'd568785526;
array[6862]=30'd839339599;
array[6863]=30'd808945195;
array[6864]=30'd503787028;
array[6865]=30'd396842530;
array[6866]=30'd724009508;
array[6867]=30'd778553911;
array[6868]=30'd556235306;
array[6869]=30'd470243883;
array[6870]=30'd941029952;
array[6871]=30'd981941808;
array[6872]=30'd981941808;
array[6873]=30'd963075636;
array[6874]=30'd963075636;
array[6875]=30'd963075636;
array[6876]=30'd963075636;
array[6877]=30'd641178184;
array[6878]=30'd336049694;
array[6879]=30'd598167087;
array[6880]=30'd681011766;
array[6881]=30'd470243883;
array[6882]=30'd256341531;
array[6883]=30'd503787028;
array[6884]=30'd681011766;
array[6885]=30'd884420162;
array[6886]=30'd963075636;
array[6887]=30'd916923947;
array[6888]=30'd793183798;
array[6889]=30'd604358258;
array[6890]=30'd634745492;
array[6891]=30'd444952244;
array[6892]=30'd608524977;
array[6893]=30'd644157123;
array[6894]=30'd581260986;
array[6895]=30'd553991871;
array[6896]=30'd644157123;
array[6897]=30'd548772504;
array[6898]=30'd852917899;
array[6899]=30'd852917899;
array[6900]=30'd852917899;
array[6901]=30'd852917899;
array[6902]=30'd852917899;
array[6903]=30'd852917899;
array[6904]=30'd852917899;
array[6905]=30'd852917899;
array[6906]=30'd852917899;
array[6907]=30'd852917899;
array[6908]=30'd852917899;
array[6909]=30'd852917899;
array[6910]=30'd852917899;
array[6911]=30'd852917899;
array[6912]=30'd852917899;
array[6913]=30'd873911932;
array[6914]=30'd873911932;
array[6915]=30'd873911932;
array[6916]=30'd873911932;
array[6917]=30'd873911932;
array[6918]=30'd873911932;
array[6919]=30'd873911932;
array[6920]=30'd873911932;
array[6921]=30'd873911932;
array[6922]=30'd900139626;
array[6923]=30'd920102487;
array[6924]=30'd936883742;
array[6925]=30'd819437027;
array[6926]=30'd842495488;
array[6927]=30'd936883742;
array[6928]=30'd875032088;
array[6929]=30'd860306981;
array[6930]=30'd884420162;
array[6931]=30'd916923947;
array[6932]=30'd884420162;
array[6933]=30'd839339599;
array[6934]=30'd884420162;
array[6935]=30'd873911932;
array[6936]=30'd873911932;
array[6937]=30'd873911932;
array[6938]=30'd873911932;
array[6939]=30'd873911932;
array[6940]=30'd873911932;
array[6941]=30'd873911932;
array[6942]=30'd873911932;
array[6943]=30'd873911932;
array[6944]=30'd873911932;
array[6945]=30'd873911932;
array[6946]=30'd873911932;
array[6947]=30'd873911932;
array[6948]=30'd873911932;
array[6949]=30'd852917899;
array[6950]=30'd852917899;
array[6951]=30'd852917899;
array[6952]=30'd625394265;
array[6953]=30'd634745492;
array[6954]=30'd644157123;
array[6955]=30'd444952244;
array[6956]=30'd666226344;
array[6957]=30'd582345342;
array[6958]=30'd839339599;
array[6959]=30'd355962430;
array[6960]=30'd598167087;
array[6961]=30'd916923947;
array[6962]=30'd963075636;
array[6963]=30'd963075636;
array[6964]=30'd963075636;
array[6965]=30'd916923947;
array[6966]=30'd963075636;
array[6967]=30'd963075636;
array[6968]=30'd963075636;
array[6969]=30'd963075636;
array[6970]=30'd963075636;
array[6971]=30'd963075636;
array[6972]=30'd963075636;
array[6973]=30'd860306981;
array[6974]=30'd916923947;
array[6975]=30'd963075636;
array[6976]=30'd963075636;
array[6977]=30'd963075636;
array[6978]=30'd808945195;
array[6979]=30'd470243883;
array[6980]=30'd316077611;
array[6981]=30'd860306981;
array[6982]=30'd963075636;
array[6983]=30'd941029952;
array[6984]=30'd756500033;
array[6985]=30'd604358258;
array[6986]=30'd608524977;
array[6987]=30'd461756049;
array[6988]=30'd516257448;
array[6989]=30'd644157123;
array[6990]=30'd525668044;
array[6991]=30'd581260986;
array[6992]=30'd608524977;
array[6993]=30'd650530435;
array[6994]=30'd884420162;
array[6995]=30'd873911932;
array[6996]=30'd873911932;
array[6997]=30'd873911932;
array[6998]=30'd873911932;
array[6999]=30'd873911932;
array[7000]=30'd873911932;
array[7001]=30'd873911932;
array[7002]=30'd873911932;
array[7003]=30'd873911932;
array[7004]=30'd852917899;
array[7005]=30'd852917899;
array[7006]=30'd852917899;
array[7007]=30'd852917899;
array[7008]=30'd852917899;
array[7009]=30'd873911932;
array[7010]=30'd873911932;
array[7011]=30'd873911932;
array[7012]=30'd873911932;
array[7013]=30'd873911932;
array[7014]=30'd873911932;
array[7015]=30'd873911932;
array[7016]=30'd873911932;
array[7017]=30'd900139626;
array[7018]=30'd920102487;
array[7019]=30'd963075636;
array[7020]=30'd896012764;
array[7021]=30'd776468978;
array[7022]=30'd884422147;
array[7023]=30'd1002945052;
array[7024]=30'd855119352;
array[7025]=30'd776468978;
array[7026]=30'd875032088;
array[7027]=30'd963077644;
array[7028]=30'd875032088;
array[7029]=30'd842495488;
array[7030]=30'd860306981;
array[7031]=30'd884420162;
array[7032]=30'd873911932;
array[7033]=30'd873911932;
array[7034]=30'd873911932;
array[7035]=30'd873911932;
array[7036]=30'd873911932;
array[7037]=30'd873911932;
array[7038]=30'd873911932;
array[7039]=30'd873911932;
array[7040]=30'd873911932;
array[7041]=30'd873911932;
array[7042]=30'd873911932;
array[7043]=30'd873911932;
array[7044]=30'd873911932;
array[7045]=30'd873911932;
array[7046]=30'd873911932;
array[7047]=30'd873911932;
array[7048]=30'd683036269;
array[7049]=30'd634745492;
array[7050]=30'd661993129;
array[7051]=30'd485848753;
array[7052]=30'd666226344;
array[7053]=30'd559296136;
array[7054]=30'd641178184;
array[7055]=30'd613919272;
array[7056]=30'd963075636;
array[7057]=30'd963075636;
array[7058]=30'd963075636;
array[7059]=30'd963075636;
array[7060]=30'd963075636;
array[7061]=30'd963075636;
array[7062]=30'd963075636;
array[7063]=30'd963075636;
array[7064]=30'd963075636;
array[7065]=30'd963075636;
array[7066]=30'd981941808;
array[7067]=30'd963075636;
array[7068]=30'd963075636;
array[7069]=30'd963075636;
array[7070]=30'd963075636;
array[7071]=30'd963075636;
array[7072]=30'd963075636;
array[7073]=30'd963075636;
array[7074]=30'd963075636;
array[7075]=30'd916923947;
array[7076]=30'd556235306;
array[7077]=30'd396842530;
array[7078]=30'd963075636;
array[7079]=30'd941029952;
array[7080]=30'd664186439;
array[7081]=30'd625322602;
array[7082]=30'd608524977;
array[7083]=30'd394645149;
array[7084]=30'd548772504;
array[7085]=30'd644157123;
array[7086]=30'd516257448;
array[7087]=30'd608524977;
array[7088]=30'd608524977;
array[7089]=30'd710361687;
array[7090]=30'd941029952;
array[7091]=30'd884420162;
array[7092]=30'd900139626;
array[7093]=30'd900139626;
array[7094]=30'd941029952;
array[7095]=30'd963075636;
array[7096]=30'd963075636;
array[7097]=30'd963075636;
array[7098]=30'd941029952;
array[7099]=30'd900139626;
array[7100]=30'd873911932;
array[7101]=30'd852917899;
array[7102]=30'd852917899;
array[7103]=30'd852917899;
array[7104]=30'd873911932;
array[7105]=30'd873911932;
array[7106]=30'd873911932;
array[7107]=30'd873911932;
array[7108]=30'd873911932;
array[7109]=30'd873911932;
array[7110]=30'd873911932;
array[7111]=30'd873911932;
array[7112]=30'd873911932;
array[7113]=30'd900139626;
array[7114]=30'd963075636;
array[7115]=30'd936883742;
array[7116]=30'd785935846;
array[7117]=30'd819437027;
array[7118]=30'd884422147;
array[7119]=30'd983039487;
array[7120]=30'd855119352;
array[7121]=30'd754446794;
array[7122]=30'd842495488;
array[7123]=30'd946320871;
array[7124]=30'd896012764;
array[7125]=30'd754446794;
array[7126]=30'd842495488;
array[7127]=30'd884420162;
array[7128]=30'd873911932;
array[7129]=30'd873911932;
array[7130]=30'd873911932;
array[7131]=30'd873911932;
array[7132]=30'd873911932;
array[7133]=30'd873911932;
array[7134]=30'd873911932;
array[7135]=30'd873911932;
array[7136]=30'd873911932;
array[7137]=30'd873911932;
array[7138]=30'd873911932;
array[7139]=30'd873911932;
array[7140]=30'd873911932;
array[7141]=30'd873911932;
array[7142]=30'd873911932;
array[7143]=30'd873911932;
array[7144]=30'd734429821;
array[7145]=30'd591795877;
array[7146]=30'd661993129;
array[7147]=30'd496374434;
array[7148]=30'd666226344;
array[7149]=30'd568785526;
array[7150]=30'd916923947;
array[7151]=30'd920102487;
array[7152]=30'd963075636;
array[7153]=30'd963075636;
array[7154]=30'd963075636;
array[7155]=30'd963075636;
array[7156]=30'd963075636;
array[7157]=30'd963075636;
array[7158]=30'd963075636;
array[7159]=30'd963075636;
array[7160]=30'd963075636;
array[7161]=30'd963075636;
array[7162]=30'd963075636;
array[7163]=30'd963075636;
array[7164]=30'd963075636;
array[7165]=30'd963075636;
array[7166]=30'd963075636;
array[7167]=30'd963075636;
array[7168]=30'd963075636;
array[7169]=30'd963075636;
array[7170]=30'd963075636;
array[7171]=30'd963075636;
array[7172]=30'd941029952;
array[7173]=30'd808945195;
array[7174]=30'd963075636;
array[7175]=30'd941029952;
array[7176]=30'd625394265;
array[7177]=30'd634745492;
array[7178]=30'd581260986;
array[7179]=30'd362128040;
array[7180]=30'd608524977;
array[7181]=30'd644157123;
array[7182]=30'd485848753;
array[7183]=30'd661993129;
array[7184]=30'd548772504;
array[7185]=30'd791076458;
array[7186]=30'd963075636;
array[7187]=30'd916923947;
array[7188]=30'd875032088;
array[7189]=30'd855119352;
array[7190]=30'd832058842;
array[7191]=30'd832058842;
array[7192]=30'd870853059;
array[7193]=30'd926409165;
array[7194]=30'd963077644;
array[7195]=30'd941029952;
array[7196]=30'd873911932;
array[7197]=30'd852917899;
array[7198]=30'd852917899;
array[7199]=30'd873911932;
array[7200]=30'd873911932;
array[7201]=30'd873911932;
array[7202]=30'd873911932;
array[7203]=30'd873911932;
array[7204]=30'd873911932;
array[7205]=30'd873911932;
array[7206]=30'd873911932;
array[7207]=30'd873911932;
array[7208]=30'd873911932;
array[7209]=30'd900139626;
array[7210]=30'd963075636;
array[7211]=30'd819475993;
array[7212]=30'd776468978;
array[7213]=30'd884422147;
array[7214]=30'd884422147;
array[7215]=30'd963077644;
array[7216]=30'd855119352;
array[7217]=30'd754446794;
array[7218]=30'd819437027;
array[7219]=30'd963077644;
array[7220]=30'd915924476;
array[7221]=30'd764966339;
array[7222]=30'd819437027;
array[7223]=30'd884420162;
array[7224]=30'd873911932;
array[7225]=30'd873911932;
array[7226]=30'd873911932;
array[7227]=30'd873911932;
array[7228]=30'd873911932;
array[7229]=30'd873911932;
array[7230]=30'd873911932;
array[7231]=30'd873911932;
array[7232]=30'd873911932;
array[7233]=30'd873911932;
array[7234]=30'd873911932;
array[7235]=30'd873911932;
array[7236]=30'd873911932;
array[7237]=30'd873911932;
array[7238]=30'd873911932;
array[7239]=30'd873911932;
array[7240]=30'd777409151;
array[7241]=30'd548772504;
array[7242]=30'd661993129;
array[7243]=30'd444952244;
array[7244]=30'd666226344;
array[7245]=30'd568785526;
array[7246]=30'd839339599;
array[7247]=30'd916923947;
array[7248]=30'd884420162;
array[7249]=30'd916923947;
array[7250]=30'd941029952;
array[7251]=30'd916923947;
array[7252]=30'd963075636;
array[7253]=30'd963075636;
array[7254]=30'd963075636;
array[7255]=30'd963075636;
array[7256]=30'd963075636;
array[7257]=30'd963075636;
array[7258]=30'd963075636;
array[7259]=30'd963075636;
array[7260]=30'd963075636;
array[7261]=30'd963075636;
array[7262]=30'd963075636;
array[7263]=30'd963075636;
array[7264]=30'd963075636;
array[7265]=30'd884420162;
array[7266]=30'd963075636;
array[7267]=30'd941029952;
array[7268]=30'd884420162;
array[7269]=30'd963075636;
array[7270]=30'd941029952;
array[7271]=30'd916923947;
array[7272]=30'd530993763;
array[7273]=30'd634745492;
array[7274]=30'd553991871;
array[7275]=30'd427157133;
array[7276]=30'd661993129;
array[7277]=30'd661993129;
array[7278]=30'd516257448;
array[7279]=30'd661993129;
array[7280]=30'd525726362;
array[7281]=30'd808945195;
array[7282]=30'd842495488;
array[7283]=30'd776468978;
array[7284]=30'd764966339;
array[7285]=30'd764966339;
array[7286]=30'd764966339;
array[7287]=30'd790145435;
array[7288]=30'd790145435;
array[7289]=30'd790145435;
array[7290]=30'd870853059;
array[7291]=30'd963077644;
array[7292]=30'd916923947;
array[7293]=30'd873911932;
array[7294]=30'd852917899;
array[7295]=30'd873911932;
array[7296]=30'd873911932;
array[7297]=30'd873911932;
array[7298]=30'd873911932;
array[7299]=30'd873911932;
array[7300]=30'd873911932;
array[7301]=30'd873911932;
array[7302]=30'd873911932;
array[7303]=30'd873911932;
array[7304]=30'd873911932;
array[7305]=30'd873911932;
array[7306]=30'd920102487;
array[7307]=30'd839339599;
array[7308]=30'd860306981;
array[7309]=30'd884420162;
array[7310]=30'd916923947;
array[7311]=30'd936883742;
array[7312]=30'd819475993;
array[7313]=30'd776468978;
array[7314]=30'd884422147;
array[7315]=30'd916923947;
array[7316]=30'd898096696;
array[7317]=30'd842495488;
array[7318]=30'd860306981;
array[7319]=30'd884420162;
array[7320]=30'd873911932;
array[7321]=30'd873911932;
array[7322]=30'd873911932;
array[7323]=30'd873911932;
array[7324]=30'd873911932;
array[7325]=30'd873911932;
array[7326]=30'd873911932;
array[7327]=30'd873911932;
array[7328]=30'd873911932;
array[7329]=30'd873911932;
array[7330]=30'd873911932;
array[7331]=30'd873911932;
array[7332]=30'd873911932;
array[7333]=30'd873911932;
array[7334]=30'd873911932;
array[7335]=30'd873911932;
array[7336]=30'd815162003;
array[7337]=30'd525726362;
array[7338]=30'd661993129;
array[7339]=30'd452327079;
array[7340]=30'd608524977;
array[7341]=30'd589750888;
array[7342]=30'd941029952;
array[7343]=30'd963075636;
array[7344]=30'd884420162;
array[7345]=30'd963075636;
array[7346]=30'd963075636;
array[7347]=30'd963075636;
array[7348]=30'd963075636;
array[7349]=30'd963075636;
array[7350]=30'd963075636;
array[7351]=30'd963075636;
array[7352]=30'd963075636;
array[7353]=30'd963075636;
array[7354]=30'd963075636;
array[7355]=30'd963075636;
array[7356]=30'd963075636;
array[7357]=30'd963075636;
array[7358]=30'd963075636;
array[7359]=30'd963075636;
array[7360]=30'd916923947;
array[7361]=30'd941029952;
array[7362]=30'd963075636;
array[7363]=30'd884420162;
array[7364]=30'd963075636;
array[7365]=30'd963075636;
array[7366]=30'd839339599;
array[7367]=30'd860306981;
array[7368]=30'd530993763;
array[7369]=30'd634745492;
array[7370]=30'd525726362;
array[7371]=30'd496374434;
array[7372]=30'd661993129;
array[7373]=30'd581260986;
array[7374]=30'd525668044;
array[7375]=30'd608524977;
array[7376]=30'd568785526;
array[7377]=30'd860306981;
array[7378]=30'd776468978;
array[7379]=30'd785935846;
array[7380]=30'd832058842;
array[7381]=30'd870853059;
array[7382]=30'd894973365;
array[7383]=30'd914919842;
array[7384]=30'd914919842;
array[7385]=30'd854099361;
array[7386]=30'd790145435;
array[7387]=30'd926409165;
array[7388]=30'd963077644;
array[7389]=30'd884420162;
array[7390]=30'd873911932;
array[7391]=30'd852917899;
array[7392]=30'd873911932;
array[7393]=30'd873911932;
array[7394]=30'd873911932;
array[7395]=30'd873911932;
array[7396]=30'd873911932;
array[7397]=30'd873911932;
array[7398]=30'd873911932;
array[7399]=30'd873911932;
array[7400]=30'd873911932;
array[7401]=30'd873911932;
array[7402]=30'd900139626;
array[7403]=30'd900139626;
array[7404]=30'd900139626;
array[7405]=30'd873911932;
array[7406]=30'd900139626;
array[7407]=30'd920102487;
array[7408]=30'd851962439;
array[7409]=30'd860306981;
array[7410]=30'd884420162;
array[7411]=30'd884420162;
array[7412]=30'd884420162;
array[7413]=30'd884420162;
array[7414]=30'd884420162;
array[7415]=30'd900139626;
array[7416]=30'd873911932;
array[7417]=30'd873911932;
array[7418]=30'd873911932;
array[7419]=30'd873911932;
array[7420]=30'd873911932;
array[7421]=30'd873911932;
array[7422]=30'd873911932;
array[7423]=30'd873911932;
array[7424]=30'd873911932;
array[7425]=30'd873911932;
array[7426]=30'd873911932;
array[7427]=30'd873911932;
array[7428]=30'd873911932;
array[7429]=30'd873911932;
array[7430]=30'd873911932;
array[7431]=30'd873911932;
array[7432]=30'd852917899;
array[7433]=30'd525726362;
array[7434]=30'd634745492;
array[7435]=30'd452327079;
array[7436]=30'd615902883;
array[7437]=30'd734429821;
array[7438]=30'd963075636;
array[7439]=30'd963075636;
array[7440]=30'd963075636;
array[7441]=30'd963075636;
array[7442]=30'd963075636;
array[7443]=30'd963075636;
array[7444]=30'd963075636;
array[7445]=30'd963075636;
array[7446]=30'd963075636;
array[7447]=30'd963075636;
array[7448]=30'd981941808;
array[7449]=30'd963075636;
array[7450]=30'd963075636;
array[7451]=30'd963075636;
array[7452]=30'd963075636;
array[7453]=30'd963075636;
array[7454]=30'd963075636;
array[7455]=30'd963075636;
array[7456]=30'd963075636;
array[7457]=30'd963075636;
array[7458]=30'd963075636;
array[7459]=30'd963075636;
array[7460]=30'd963075636;
array[7461]=30'd963075636;
array[7462]=30'd941029952;
array[7463]=30'd793183798;
array[7464]=30'd582345342;
array[7465]=30'd634745492;
array[7466]=30'd461756049;
array[7467]=30'd553991871;
array[7468]=30'd661993129;
array[7469]=30'd516257448;
array[7470]=30'd615902883;
array[7471]=30'd615902883;
array[7472]=30'd641178184;
array[7473]=30'd819475993;
array[7474]=30'd764966339;
array[7475]=30'd894973365;
array[7476]=30'd855119352;
array[7477]=30'd832058842;
array[7478]=30'd810051001;
array[7479]=30'd778588583;
array[7480]=30'd790145435;
array[7481]=30'd834187654;
array[7482]=30'd790145435;
array[7483]=30'd870853059;
array[7484]=30'd963077644;
array[7485]=30'd884420162;
array[7486]=30'd873911932;
array[7487]=30'd873911932;
array[7488]=30'd900139626;
array[7489]=30'd873911932;
array[7490]=30'd873911932;
array[7491]=30'd873911932;
array[7492]=30'd873911932;
array[7493]=30'd873911932;
array[7494]=30'd873911932;
array[7495]=30'd900139626;
array[7496]=30'd873911932;
array[7497]=30'd873911932;
array[7498]=30'd873911932;
array[7499]=30'd900139626;
array[7500]=30'd900139626;
array[7501]=30'd900139626;
array[7502]=30'd900139626;
array[7503]=30'd900139626;
array[7504]=30'd900139626;
array[7505]=30'd873911932;
array[7506]=30'd900139626;
array[7507]=30'd873911932;
array[7508]=30'd873911932;
array[7509]=30'd900139626;
array[7510]=30'd900139626;
array[7511]=30'd873911932;
array[7512]=30'd873911932;
array[7513]=30'd873911932;
array[7514]=30'd873911932;
array[7515]=30'd873911932;
array[7516]=30'd873911932;
array[7517]=30'd873911932;
array[7518]=30'd873911932;
array[7519]=30'd873911932;
array[7520]=30'd873911932;
array[7521]=30'd873911932;
array[7522]=30'd873911932;
array[7523]=30'd873911932;
array[7524]=30'd873911932;
array[7525]=30'd873911932;
array[7526]=30'd873911932;
array[7527]=30'd873911932;
array[7528]=30'd873911932;
array[7529]=30'd604358258;
array[7530]=30'd634745492;
array[7531]=30'd452327079;
array[7532]=30'd591795877;
array[7533]=30'd820432476;
array[7534]=30'd963075636;
array[7535]=30'd963075636;
array[7536]=30'd963075636;
array[7537]=30'd963075636;
array[7538]=30'd963075636;
array[7539]=30'd963075636;
array[7540]=30'd963075636;
array[7541]=30'd963075636;
array[7542]=30'd963075636;
array[7543]=30'd963075636;
array[7544]=30'd963075636;
array[7545]=30'd963075636;
array[7546]=30'd963075636;
array[7547]=30'd963075636;
array[7548]=30'd963075636;
array[7549]=30'd963075636;
array[7550]=30'd963075636;
array[7551]=30'd963075636;
array[7552]=30'd963075636;
array[7553]=30'd963075636;
array[7554]=30'd963075636;
array[7555]=30'd963075636;
array[7556]=30'd963075636;
array[7557]=30'd941029952;
array[7558]=30'd941029952;
array[7559]=30'd739680847;
array[7560]=30'd604358258;
array[7561]=30'd608524977;
array[7562]=30'd461756049;
array[7563]=30'd608524977;
array[7564]=30'd608524977;
array[7565]=30'd461756049;
array[7566]=30'd608524977;
array[7567]=30'd582345342;
array[7568]=30'd710361687;
array[7569]=30'd785935846;
array[7570]=30'd832058842;
array[7571]=30'd926409165;
array[7572]=30'd832058842;
array[7573]=30'd764966339;
array[7574]=30'd810051001;
array[7575]=30'd790145435;
array[7576]=30'd763929993;
array[7577]=30'd790145435;
array[7578]=30'd854099361;
array[7579]=30'd790145435;
array[7580]=30'd946320871;
array[7581]=30'd916923947;
array[7582]=30'd884420162;
array[7583]=30'd873911932;
array[7584]=30'd884420162;
array[7585]=30'd860306981;
array[7586]=30'd884420162;
array[7587]=30'd884420162;
array[7588]=30'd900139626;
array[7589]=30'd900139626;
array[7590]=30'd873911932;
array[7591]=30'd873911932;
array[7592]=30'd900139626;
array[7593]=30'd900139626;
array[7594]=30'd873911932;
array[7595]=30'd900139626;
array[7596]=30'd873911932;
array[7597]=30'd900139626;
array[7598]=30'd900139626;
array[7599]=30'd900139626;
array[7600]=30'd873911932;
array[7601]=30'd873911932;
array[7602]=30'd900139626;
array[7603]=30'd873911932;
array[7604]=30'd873911932;
array[7605]=30'd900139626;
array[7606]=30'd900139626;
array[7607]=30'd873911932;
array[7608]=30'd873911932;
array[7609]=30'd873911932;
array[7610]=30'd873911932;
array[7611]=30'd900139626;
array[7612]=30'd873911932;
array[7613]=30'd873911932;
array[7614]=30'd900139626;
array[7615]=30'd873911932;
array[7616]=30'd873911932;
array[7617]=30'd873911932;
array[7618]=30'd900139626;
array[7619]=30'd873911932;
array[7620]=30'd873911932;
array[7621]=30'd873911932;
array[7622]=30'd873911932;
array[7623]=30'd873911932;
array[7624]=30'd873911932;
array[7625]=30'd702982791;
array[7626]=30'd582345342;
array[7627]=30'd461756049;
array[7628]=30'd591795877;
array[7629]=30'd820432476;
array[7630]=30'd963075636;
array[7631]=30'd963075636;
array[7632]=30'd963075636;
array[7633]=30'd963075636;
array[7634]=30'd963075636;
array[7635]=30'd963075636;
array[7636]=30'd941029952;
array[7637]=30'd860306981;
array[7638]=30'd916923947;
array[7639]=30'd941029952;
array[7640]=30'd963075636;
array[7641]=30'd963075636;
array[7642]=30'd963075636;
array[7643]=30'd963075636;
array[7644]=30'd963075636;
array[7645]=30'd916923947;
array[7646]=30'd860306981;
array[7647]=30'd963075636;
array[7648]=30'd963075636;
array[7649]=30'd963075636;
array[7650]=30'd963075636;
array[7651]=30'd963075636;
array[7652]=30'd963075636;
array[7653]=30'd941029952;
array[7654]=30'd941029952;
array[7655]=30'd625394265;
array[7656]=30'd634745492;
array[7657]=30'd634745492;
array[7658]=30'd525726362;
array[7659]=30'd608524977;
array[7660]=30'd548772504;
array[7661]=30'd461756049;
array[7662]=30'd634745492;
array[7663]=30'd559296136;
array[7664]=30'd808945195;
array[7665]=30'd764966339;
array[7666]=30'd894973365;
array[7667]=30'd896012764;
array[7668]=30'd832058842;
array[7669]=30'd764966339;
array[7670]=30'd944268729;
array[7671]=30'd944268729;
array[7672]=30'd810051001;
array[7673]=30'd790145435;
array[7674]=30'd914919842;
array[7675]=30'd790145435;
array[7676]=30'd870853059;
array[7677]=30'd963077644;
array[7678]=30'd884420162;
array[7679]=30'd873911932;
array[7680]=30'd842495488;
array[7681]=30'd884422147;
array[7682]=30'd884422147;
array[7683]=30'd884422147;
array[7684]=30'd884420162;
array[7685]=30'd900139626;
array[7686]=30'd873911932;
array[7687]=30'd873911932;
array[7688]=30'd900139626;
array[7689]=30'd873911932;
array[7690]=30'd873911932;
array[7691]=30'd873911932;
array[7692]=30'd873911932;
array[7693]=30'd900139626;
array[7694]=30'd900139626;
array[7695]=30'd900139626;
array[7696]=30'd900139626;
array[7697]=30'd900139626;
array[7698]=30'd900139626;
array[7699]=30'd900139626;
array[7700]=30'd900139626;
array[7701]=30'd873911932;
array[7702]=30'd900139626;
array[7703]=30'd900139626;
array[7704]=30'd900139626;
array[7705]=30'd900139626;
array[7706]=30'd873911932;
array[7707]=30'd900139626;
array[7708]=30'd873911932;
array[7709]=30'd900139626;
array[7710]=30'd900139626;
array[7711]=30'd873911932;
array[7712]=30'd873911932;
array[7713]=30'd873911932;
array[7714]=30'd873911932;
array[7715]=30'd900139626;
array[7716]=30'd900139626;
array[7717]=30'd873911932;
array[7718]=30'd873911932;
array[7719]=30'd873911932;
array[7720]=30'd873911932;
array[7721]=30'd777409151;
array[7722]=30'd530993763;
array[7723]=30'd461756049;
array[7724]=30'd666226344;
array[7725]=30'd683036269;
array[7726]=30'd963075636;
array[7727]=30'd963075636;
array[7728]=30'd963075636;
array[7729]=30'd963075636;
array[7730]=30'd963075636;
array[7731]=30'd963075636;
array[7732]=30'd963075636;
array[7733]=30'd916923947;
array[7734]=30'd860306981;
array[7735]=30'd793183798;
array[7736]=30'd793183798;
array[7737]=30'd793183798;
array[7738]=30'd808945195;
array[7739]=30'd793183798;
array[7740]=30'd756500033;
array[7741]=30'd808945195;
array[7742]=30'd916923947;
array[7743]=30'd963075636;
array[7744]=30'd963075636;
array[7745]=30'd963075636;
array[7746]=30'd981941808;
array[7747]=30'd963075636;
array[7748]=30'd963075636;
array[7749]=30'd963075636;
array[7750]=30'd916923947;
array[7751]=30'd556154453;
array[7752]=30'd665151100;
array[7753]=30'd548772504;
array[7754]=30'd608524977;
array[7755]=30'd608524977;
array[7756]=30'd427157133;
array[7757]=30'd525726362;
array[7758]=30'd634745492;
array[7759]=30'd559296136;
array[7760]=30'd819475993;
array[7761]=30'd810051001;
array[7762]=30'd926409165;
array[7763]=30'd884422147;
array[7764]=30'd819475993;
array[7765]=30'd764966339;
array[7766]=30'd944268729;
array[7767]=30'd894973365;
array[7768]=30'd810051001;
array[7769]=30'd790145435;
array[7770]=30'd914919842;
array[7771]=30'd790145435;
array[7772]=30'd870853059;
array[7773]=30'd915924476;
array[7774]=30'd884420162;
array[7775]=30'd873911932;
array[7776]=30'd870853059;
array[7777]=30'd896012764;
array[7778]=30'd855119352;
array[7779]=30'd884422147;
array[7780]=30'd884420162;
array[7781]=30'd900139626;
array[7782]=30'd900139626;
array[7783]=30'd900139626;
array[7784]=30'd873911932;
array[7785]=30'd873911932;
array[7786]=30'd873911932;
array[7787]=30'd873911932;
array[7788]=30'd873911932;
array[7789]=30'd900139626;
array[7790]=30'd900139626;
array[7791]=30'd900139626;
array[7792]=30'd900139626;
array[7793]=30'd900139626;
array[7794]=30'd900139626;
array[7795]=30'd900139626;
array[7796]=30'd900139626;
array[7797]=30'd900139626;
array[7798]=30'd900139626;
array[7799]=30'd900139626;
array[7800]=30'd900139626;
array[7801]=30'd900139626;
array[7802]=30'd900139626;
array[7803]=30'd900139626;
array[7804]=30'd900139626;
array[7805]=30'd900139626;
array[7806]=30'd900139626;
array[7807]=30'd873911932;
array[7808]=30'd873911932;
array[7809]=30'd900139626;
array[7810]=30'd900139626;
array[7811]=30'd900139626;
array[7812]=30'd900139626;
array[7813]=30'd873911932;
array[7814]=30'd873911932;
array[7815]=30'd873911932;
array[7816]=30'd873911932;
array[7817]=30'd873911932;
array[7818]=30'd503733877;
array[7819]=30'd484819572;
array[7820]=30'd661993129;
array[7821]=30'd591795877;
array[7822]=30'd820432476;
array[7823]=30'd963075636;
array[7824]=30'd963075636;
array[7825]=30'd963075636;
array[7826]=30'd963075636;
array[7827]=30'd963075636;
array[7828]=30'd963075636;
array[7829]=30'd963075636;
array[7830]=30'd963075636;
array[7831]=30'd963075636;
array[7832]=30'd981941808;
array[7833]=30'd981941808;
array[7834]=30'd981941808;
array[7835]=30'd963075636;
array[7836]=30'd963075636;
array[7837]=30'd963075636;
array[7838]=30'd963075636;
array[7839]=30'd963075636;
array[7840]=30'd963075636;
array[7841]=30'd963075636;
array[7842]=30'd963075636;
array[7843]=30'd963075636;
array[7844]=30'd963075636;
array[7845]=30'd941029952;
array[7846]=30'd884420162;
array[7847]=30'd530993763;
array[7848]=30'd634745492;
array[7849]=30'd444952244;
array[7850]=30'd661993129;
array[7851]=30'd553991871;
array[7852]=30'd331722417;
array[7853]=30'd591795877;
array[7854]=30'd615902883;
array[7855]=30'd589750888;
array[7856]=30'd819475993;
array[7857]=30'd810051001;
array[7858]=30'd946320871;
array[7859]=30'd875032088;
array[7860]=30'd819475993;
array[7861]=30'd764966339;
array[7862]=30'd894973365;
array[7863]=30'd810051001;
array[7864]=30'd764966339;
array[7865]=30'd778588583;
array[7866]=30'd883468684;
array[7867]=30'd790145435;
array[7868]=30'd870853059;
array[7869]=30'd915924476;
array[7870]=30'd884420162;
array[7871]=30'd873911932;
array[7872]=30'd855119352;
array[7873]=30'd855119352;
array[7874]=30'd884422147;
array[7875]=30'd916923947;
array[7876]=30'd884420162;
array[7877]=30'd900139626;
array[7878]=30'd900139626;
array[7879]=30'd900139626;
array[7880]=30'd900139626;
array[7881]=30'd900139626;
array[7882]=30'd900139626;
array[7883]=30'd900139626;
array[7884]=30'd900139626;
array[7885]=30'd900139626;
array[7886]=30'd900139626;
array[7887]=30'd900139626;
array[7888]=30'd900139626;
array[7889]=30'd900139626;
array[7890]=30'd900139626;
array[7891]=30'd900139626;
array[7892]=30'd900139626;
array[7893]=30'd900139626;
array[7894]=30'd900139626;
array[7895]=30'd900139626;
array[7896]=30'd900139626;
array[7897]=30'd900139626;
array[7898]=30'd900139626;
array[7899]=30'd900139626;
array[7900]=30'd900139626;
array[7901]=30'd900139626;
array[7902]=30'd900139626;
array[7903]=30'd900139626;
array[7904]=30'd900139626;
array[7905]=30'd900139626;
array[7906]=30'd900139626;
array[7907]=30'd900139626;
array[7908]=30'd900139626;
array[7909]=30'd873911932;
array[7910]=30'd873911932;
array[7911]=30'd873911932;
array[7912]=30'd873911932;
array[7913]=30'd873911932;
array[7914]=30'd530993763;
array[7915]=30'd447089265;
array[7916]=30'd661993129;
array[7917]=30'd608524977;
array[7918]=30'd433483392;
array[7919]=30'd739680847;
array[7920]=30'd941029952;
array[7921]=30'd963075636;
array[7922]=30'd963075636;
array[7923]=30'd963075636;
array[7924]=30'd963075636;
array[7925]=30'd963075636;
array[7926]=30'd963075636;
array[7927]=30'd963075636;
array[7928]=30'd963075636;
array[7929]=30'd981941808;
array[7930]=30'd963075636;
array[7931]=30'd963075636;
array[7932]=30'd963075636;
array[7933]=30'd963075636;
array[7934]=30'd963075636;
array[7935]=30'd963075636;
array[7936]=30'd963075636;
array[7937]=30'd963075636;
array[7938]=30'd963075636;
array[7939]=30'd963075636;
array[7940]=30'd963075636;
array[7941]=30'd941029952;
array[7942]=30'd625394265;
array[7943]=30'd582345342;
array[7944]=30'd548772504;
array[7945]=30'd553991871;
array[7946]=30'd608524977;
array[7947]=30'd452327079;
array[7948]=30'd394645149;
array[7949]=30'd634745492;
array[7950]=30'd591795877;
array[7951]=30'd674710128;
array[7952]=30'd819475993;
array[7953]=30'd810051001;
array[7954]=30'd963129822;
array[7955]=30'd936883742;
array[7956]=30'd855119352;
array[7957]=30'd764966339;
array[7958]=30'd894973365;
array[7959]=30'd944268729;
array[7960]=30'd870853059;
array[7961]=30'd854099361;
array[7962]=30'd790145435;
array[7963]=30'd778588583;
array[7964]=30'd896012764;
array[7965]=30'd884422147;
array[7966]=30'd873911932;
array[7967]=30'd873911932;
array[7968]=30'd875032088;
array[7969]=30'd884422147;
array[7970]=30'd884422147;
array[7971]=30'd884420162;
array[7972]=30'd900139626;
array[7973]=30'd900139626;
array[7974]=30'd900139626;
array[7975]=30'd900139626;
array[7976]=30'd900139626;
array[7977]=30'd900139626;
array[7978]=30'd900139626;
array[7979]=30'd900139626;
array[7980]=30'd900139626;
array[7981]=30'd900139626;
array[7982]=30'd900139626;
array[7983]=30'd900139626;
array[7984]=30'd900139626;
array[7985]=30'd900139626;
array[7986]=30'd900139626;
array[7987]=30'd900139626;
array[7988]=30'd900139626;
array[7989]=30'd900139626;
array[7990]=30'd900139626;
array[7991]=30'd900139626;
array[7992]=30'd900139626;
array[7993]=30'd900139626;
array[7994]=30'd900139626;
array[7995]=30'd900139626;
array[7996]=30'd900139626;
array[7997]=30'd900139626;
array[7998]=30'd900139626;
array[7999]=30'd900139626;
array[8000]=30'd900139626;
array[8001]=30'd900139626;
array[8002]=30'd900139626;
array[8003]=30'd900139626;
array[8004]=30'd900139626;
array[8005]=30'd900139626;
array[8006]=30'd900139626;
array[8007]=30'd873911932;
array[8008]=30'd873911932;
array[8009]=30'd873911932;
array[8010]=30'd625394265;
array[8011]=30'd447089265;
array[8012]=30'd661993129;
array[8013]=30'd608524977;
array[8014]=30'd452327079;
array[8015]=30'd433483392;
array[8016]=30'd641178184;
array[8017]=30'd884420162;
array[8018]=30'd963075636;
array[8019]=30'd963075636;
array[8020]=30'd963075636;
array[8021]=30'd963075636;
array[8022]=30'd963075636;
array[8023]=30'd963075636;
array[8024]=30'd963075636;
array[8025]=30'd981941808;
array[8026]=30'd963075636;
array[8027]=30'd963075636;
array[8028]=30'd963075636;
array[8029]=30'd963075636;
array[8030]=30'd963075636;
array[8031]=30'd963075636;
array[8032]=30'd963075636;
array[8033]=30'd963075636;
array[8034]=30'd963075636;
array[8035]=30'd963075636;
array[8036]=30'd884420162;
array[8037]=30'd625394265;
array[8038]=30'd374749802;
array[8039]=30'd634745492;
array[8040]=30'd452327079;
array[8041]=30'd608524977;
array[8042]=30'd548772504;
array[8043]=30'd331722417;
array[8044]=30'd461756049;
array[8045]=30'd634745492;
array[8046]=30'd582345342;
array[8047]=30'd744992360;
array[8048]=30'd808945195;
array[8049]=30'd785935846;
array[8050]=30'd963129822;
array[8051]=30'd983039487;
array[8052]=30'd875032088;
array[8053]=30'd764966339;
array[8054]=30'd810051001;
array[8055]=30'd944268729;
array[8056]=30'd997736898;
array[8057]=30'd944268729;
array[8058]=30'd778588583;
array[8059]=30'd810051001;
array[8060]=30'd915924476;
array[8061]=30'd884420162;
array[8062]=30'd873911932;
array[8063]=30'd873911932;
array[8064]=30'd898096696;
array[8065]=30'd884420162;
array[8066]=30'd884420162;
array[8067]=30'd884420162;
array[8068]=30'd900139626;
array[8069]=30'd900139626;
array[8070]=30'd900139626;
array[8071]=30'd900139626;
array[8072]=30'd900139626;
array[8073]=30'd900139626;
array[8074]=30'd900139626;
array[8075]=30'd900139626;
array[8076]=30'd900139626;
array[8077]=30'd900139626;
array[8078]=30'd900139626;
array[8079]=30'd900139626;
array[8080]=30'd900139626;
array[8081]=30'd900139626;
array[8082]=30'd900139626;
array[8083]=30'd900139626;
array[8084]=30'd900139626;
array[8085]=30'd900139626;
array[8086]=30'd900139626;
array[8087]=30'd900139626;
array[8088]=30'd900139626;
array[8089]=30'd900139626;
array[8090]=30'd900139626;
array[8091]=30'd900139626;
array[8092]=30'd900139626;
array[8093]=30'd900139626;
array[8094]=30'd900139626;
array[8095]=30'd900139626;
array[8096]=30'd884420162;
array[8097]=30'd884420162;
array[8098]=30'd884420162;
array[8099]=30'd884420162;
array[8100]=30'd884420162;
array[8101]=30'd900139626;
array[8102]=30'd900139626;
array[8103]=30'd873911932;
array[8104]=30'd900139626;
array[8105]=30'd873911932;
array[8106]=30'd674710128;
array[8107]=30'd484819572;
array[8108]=30'd634745492;
array[8109]=30'd553991871;
array[8110]=30'd452327079;
array[8111]=30'd427157133;
array[8112]=30'd351684214;
array[8113]=30'd456562280;
array[8114]=30'd710361687;
array[8115]=30'd916923947;
array[8116]=30'd941029952;
array[8117]=30'd963075636;
array[8118]=30'd963075636;
array[8119]=30'd963075636;
array[8120]=30'd963075636;
array[8121]=30'd963075636;
array[8122]=30'd963075636;
array[8123]=30'd963075636;
array[8124]=30'd963075636;
array[8125]=30'd963075636;
array[8126]=30'd963075636;
array[8127]=30'd963075636;
array[8128]=30'd963075636;
array[8129]=30'd963075636;
array[8130]=30'd941029952;
array[8131]=30'd756500033;
array[8132]=30'd450262593;
array[8133]=30'd421932631;
array[8134]=30'd447089265;
array[8135]=30'd582345342;
array[8136]=30'd516257448;
array[8137]=30'd581260986;
array[8138]=30'd427157133;
array[8139]=30'd328601227;
array[8140]=30'd461756049;
array[8141]=30'd634745492;
array[8142]=30'd525726362;
array[8143]=30'd839339599;
array[8144]=30'd851962439;
array[8145]=30'd785935846;
array[8146]=30'd832058842;
array[8147]=30'd963129822;
array[8148]=30'd983039487;
array[8149]=30'd832058842;
array[8150]=30'd764966339;
array[8151]=30'd764966339;
array[8152]=30'd810051001;
array[8153]=30'd778588583;
array[8154]=30'd778588583;
array[8155]=30'd896012764;
array[8156]=30'd884422147;
array[8157]=30'd884420162;
array[8158]=30'd900139626;
array[8159]=30'd873911932;
array[8160]=30'd900139626;
array[8161]=30'd884420162;
array[8162]=30'd900139626;
array[8163]=30'd900139626;
array[8164]=30'd900139626;
array[8165]=30'd900139626;
array[8166]=30'd900139626;
array[8167]=30'd900139626;
array[8168]=30'd900139626;
array[8169]=30'd900139626;
array[8170]=30'd900139626;
array[8171]=30'd900139626;
array[8172]=30'd900139626;
array[8173]=30'd900139626;
array[8174]=30'd900139626;
array[8175]=30'd900139626;
array[8176]=30'd900139626;
array[8177]=30'd900139626;
array[8178]=30'd900139626;
array[8179]=30'd900139626;
array[8180]=30'd900139626;
array[8181]=30'd900139626;
array[8182]=30'd900139626;
array[8183]=30'd900139626;
array[8184]=30'd900139626;
array[8185]=30'd900139626;
array[8186]=30'd900139626;
array[8187]=30'd900139626;
array[8188]=30'd900139626;
array[8189]=30'd900139626;
array[8190]=30'd900139626;
array[8191]=30'd900139626;
array[8192]=30'd808945195;
array[8193]=30'd936883742;
array[8194]=30'd916923947;
array[8195]=30'd819475993;
array[8196]=30'd936883742;
array[8197]=30'd941029952;
array[8198]=30'd900139626;
array[8199]=30'd900139626;
array[8200]=30'd900139626;
array[8201]=30'd873911932;
array[8202]=30'd739680847;
array[8203]=30'd530993763;
array[8204]=30'd634745492;
array[8205]=30'd553991871;
array[8206]=30'd452327079;
array[8207]=30'd461756049;
array[8208]=30'd351684214;
array[8209]=30'd456562280;
array[8210]=30'd421932631;
array[8211]=30'd421987917;
array[8212]=30'd625394265;
array[8213]=30'd793183798;
array[8214]=30'd916923947;
array[8215]=30'd941029952;
array[8216]=30'd963075636;
array[8217]=30'd963075636;
array[8218]=30'd963075636;
array[8219]=30'd963075636;
array[8220]=30'd963075636;
array[8221]=30'd963075636;
array[8222]=30'd963075636;
array[8223]=30'd963075636;
array[8224]=30'd884420162;
array[8225]=30'd756500033;
array[8226]=30'd512140869;
array[8227]=30'd450262593;
array[8228]=30'd421932631;
array[8229]=30'd397823583;
array[8230]=30'd503733877;
array[8231]=30'd461756049;
array[8232]=30'd591795877;
array[8233]=30'd496374434;
array[8234]=30'd300284569;
array[8235]=30'd260455061;
array[8236]=30'd503733877;
array[8237]=30'd634745492;
array[8238]=30'd559296136;
array[8239]=30'd873911932;
array[8240]=30'd898096696;
array[8241]=30'd819475993;
array[8242]=30'd785935846;
array[8243]=30'd896012764;
array[8244]=30'd1016593896;
array[8245]=30'd915924476;
array[8246]=30'd855119352;
array[8247]=30'd832058842;
array[8248]=30'd785935846;
array[8249]=30'd819437027;
array[8250]=30'd855119352;
array[8251]=30'd884422147;
array[8252]=30'd884420162;
array[8253]=30'd900139626;
array[8254]=30'd900139626;
array[8255]=30'd873911932;
array[8256]=30'd900139626;
array[8257]=30'd900139626;
array[8258]=30'd900139626;
array[8259]=30'd900139626;
array[8260]=30'd900139626;
array[8261]=30'd900139626;
array[8262]=30'd900139626;
array[8263]=30'd900139626;
array[8264]=30'd900139626;
array[8265]=30'd900139626;
array[8266]=30'd900139626;
array[8267]=30'd900139626;
array[8268]=30'd900139626;
array[8269]=30'd900139626;
array[8270]=30'd900139626;
array[8271]=30'd900139626;
array[8272]=30'd900139626;
array[8273]=30'd900139626;
array[8274]=30'd900139626;
array[8275]=30'd900139626;
array[8276]=30'd900139626;
array[8277]=30'd900139626;
array[8278]=30'd900139626;
array[8279]=30'd900139626;
array[8280]=30'd900139626;
array[8281]=30'd900139626;
array[8282]=30'd900139626;
array[8283]=30'd900139626;
array[8284]=30'd900139626;
array[8285]=30'd900139626;
array[8286]=30'd900139626;
array[8287]=30'd920102487;
array[8288]=30'd851962439;
array[8289]=30'd936883742;
array[8290]=30'd915924476;
array[8291]=30'd776468978;
array[8292]=30'd983039487;
array[8293]=30'd936883742;
array[8294]=30'd860306981;
array[8295]=30'd860306981;
array[8296]=30'd884420162;
array[8297]=30'd900139626;
array[8298]=30'd791076458;
array[8299]=30'd559296136;
array[8300]=30'd634745492;
array[8301]=30'd516257448;
array[8302]=30'd452327079;
array[8303]=30'd433483392;
array[8304]=30'd368466587;
array[8305]=30'd433483392;
array[8306]=30'd409379461;
array[8307]=30'd397823583;
array[8308]=30'd456562280;
array[8309]=30'd397823583;
array[8310]=30'd421987917;
array[8311]=30'd547846737;
array[8312]=30'd664186439;
array[8313]=30'd793183798;
array[8314]=30'd839339599;
array[8315]=30'd884420162;
array[8316]=30'd839339599;
array[8317]=30'd793183798;
array[8318]=30'd710361687;
array[8319]=30'd664186439;
array[8320]=30'd681011766;
array[8321]=30'd756500033;
array[8322]=30'd335980112;
array[8323]=30'd450262593;
array[8324]=30'd456562280;
array[8325]=30'd374749802;
array[8326]=30'd525726362;
array[8327]=30'd496374434;
array[8328]=30'd548772504;
array[8329]=30'd368466587;
array[8330]=30'd300284569;
array[8331]=30'd300284569;
array[8332]=30'd496374434;
array[8333]=30'd608524977;
array[8334]=30'd582345342;
array[8335]=30'd900139626;
array[8336]=30'd900139626;
array[8337]=30'd898096696;
array[8338]=30'd819475993;
array[8339]=30'd785935846;
array[8340]=30'd946320871;
array[8341]=30'd983039487;
array[8342]=30'd936883742;
array[8343]=30'd915924476;
array[8344]=30'd915924476;
array[8345]=30'd936883742;
array[8346]=30'd916923947;
array[8347]=30'd884420162;
array[8348]=30'd900139626;
array[8349]=30'd900139626;
array[8350]=30'd873911932;
array[8351]=30'd873911932;
array[8352]=30'd900139626;
array[8353]=30'd900139626;
array[8354]=30'd900139626;
array[8355]=30'd900139626;
array[8356]=30'd900139626;
array[8357]=30'd900139626;
array[8358]=30'd900139626;
array[8359]=30'd898096696;
array[8360]=30'd851962439;
array[8361]=30'd860306981;
array[8362]=30'd860306981;
array[8363]=30'd898096696;
array[8364]=30'd884420162;
array[8365]=30'd900139626;
array[8366]=30'd900139626;
array[8367]=30'd900139626;
array[8368]=30'd900139626;
array[8369]=30'd900139626;
array[8370]=30'd900139626;
array[8371]=30'd900139626;
array[8372]=30'd900139626;
array[8373]=30'd900139626;
array[8374]=30'd900139626;
array[8375]=30'd900139626;
array[8376]=30'd900139626;
array[8377]=30'd900139626;
array[8378]=30'd900139626;
array[8379]=30'd900139626;
array[8380]=30'd900139626;
array[8381]=30'd900139626;
array[8382]=30'd900139626;
array[8383]=30'd920102487;
array[8384]=30'd898096696;
array[8385]=30'd936883742;
array[8386]=30'd898096696;
array[8387]=30'd855119352;
array[8388]=30'd983039487;
array[8389]=30'd875032088;
array[8390]=30'd842495488;
array[8391]=30'd936883742;
array[8392]=30'd916923947;
array[8393]=30'd900139626;
array[8394]=30'd777409151;
array[8395]=30'd582345342;
array[8396]=30'd608524977;
array[8397]=30'd485848753;
array[8398]=30'd461756049;
array[8399]=30'd397823583;
array[8400]=30'd409379461;
array[8401]=30'd427157133;
array[8402]=30'd409379461;
array[8403]=30'd351684214;
array[8404]=30'd447089265;
array[8405]=30'd433483392;
array[8406]=30'd433483392;
array[8407]=30'd447089265;
array[8408]=30'd397823583;
array[8409]=30'd450262593;
array[8410]=30'd756500033;
array[8411]=30'd793183798;
array[8412]=30'd793183798;
array[8413]=30'd791076458;
array[8414]=30'd791076458;
array[8415]=30'd820432476;
array[8416]=30'd820432476;
array[8417]=30'd756500033;
array[8418]=30'd247985748;
array[8419]=30'd312961612;
array[8420]=30'd421932631;
array[8421]=30'd447089265;
array[8422]=30'd461756049;
array[8423]=30'd591795877;
array[8424]=30'd452327079;
array[8425]=30'd260455061;
array[8426]=30'd368466587;
array[8427]=30'd351684214;
array[8428]=30'd525726362;
array[8429]=30'd608524977;
array[8430]=30'd625394265;
array[8431]=30'd900139626;
array[8432]=30'd900139626;
array[8433]=30'd884420162;
array[8434]=30'd851962439;
array[8435]=30'd785935846;
array[8436]=30'd832058842;
array[8437]=30'd963129822;
array[8438]=30'd963129822;
array[8439]=30'd963129822;
array[8440]=30'd946320871;
array[8441]=30'd946320871;
array[8442]=30'd963075636;
array[8443]=30'd900139626;
array[8444]=30'd900139626;
array[8445]=30'd900139626;
array[8446]=30'd900139626;
array[8447]=30'd900139626;
array[8448]=30'd900139626;
array[8449]=30'd900139626;
array[8450]=30'd900139626;
array[8451]=30'd900139626;
array[8452]=30'd900139626;
array[8453]=30'd900139626;
array[8454]=30'd851962439;
array[8455]=30'd819475993;
array[8456]=30'd832058842;
array[8457]=30'd832058842;
array[8458]=30'd832058842;
array[8459]=30'd776468978;
array[8460]=30'd842495488;
array[8461]=30'd916923947;
array[8462]=30'd900139626;
array[8463]=30'd900139626;
array[8464]=30'd900139626;
array[8465]=30'd900139626;
array[8466]=30'd900139626;
array[8467]=30'd900139626;
array[8468]=30'd900139626;
array[8469]=30'd900139626;
array[8470]=30'd900139626;
array[8471]=30'd900139626;
array[8472]=30'd900139626;
array[8473]=30'd900139626;
array[8474]=30'd900139626;
array[8475]=30'd900139626;
array[8476]=30'd900139626;
array[8477]=30'd900139626;
array[8478]=30'd900139626;
array[8479]=30'd920102487;
array[8480]=30'd898096696;
array[8481]=30'd898096696;
array[8482]=30'd875032088;
array[8483]=30'd875032088;
array[8484]=30'd915924476;
array[8485]=30'd855119352;
array[8486]=30'd915924476;
array[8487]=30'd963077644;
array[8488]=30'd884420162;
array[8489]=30'd900139626;
array[8490]=30'd702982791;
array[8491]=30'd634745492;
array[8492]=30'd608524977;
array[8493]=30'd444952244;
array[8494]=30'd427157133;
array[8495]=30'd351684214;
array[8496]=30'd397823583;
array[8497]=30'd447089265;
array[8498]=30'd397823583;
array[8499]=30'd277255789;
array[8500]=30'd447089265;
array[8501]=30'd427157133;
array[8502]=30'd461756049;
array[8503]=30'd433483392;
array[8504]=30'd333912689;
array[8505]=30'd355962430;
array[8506]=30'd820432476;
array[8507]=30'd820432476;
array[8508]=30'd820432476;
array[8509]=30'd820432476;
array[8510]=30'd820432476;
array[8511]=30'd820432476;
array[8512]=30'd681011766;
array[8513]=30'd421987917;
array[8514]=30'd274187850;
array[8515]=30'd274187850;
array[8516]=30'd258398808;
array[8517]=30'd447089265;
array[8518]=30'd525726362;
array[8519]=30'd516257448;
array[8520]=30'd409379461;
array[8521]=30'd333912689;
array[8522]=30'd421932631;
array[8523]=30'd374749802;
array[8524]=30'd525726362;
array[8525]=30'd591795877;
array[8526]=30'd683036269;
array[8527]=30'd900139626;
array[8528]=30'd900139626;
array[8529]=30'd900139626;
array[8530]=30'd920102487;
array[8531]=30'd875032088;
array[8532]=30'd776468978;
array[8533]=30'd764966339;
array[8534]=30'd778588583;
array[8535]=30'd778588583;
array[8536]=30'd794287561;
array[8537]=30'd819437027;
array[8538]=30'd916923947;
array[8539]=30'd900139626;
array[8540]=30'd900139626;
array[8541]=30'd873911932;
array[8542]=30'd873911932;
array[8543]=30'd873911932;
array[8544]=30'd900139626;
array[8545]=30'd900139626;
array[8546]=30'd900139626;
array[8547]=30'd900139626;
array[8548]=30'd900139626;
array[8549]=30'd900139626;
array[8550]=30'd936883742;
array[8551]=30'd936883742;
array[8552]=30'd983039487;
array[8553]=30'd983039487;
array[8554]=30'd983039487;
array[8555]=30'd915924476;
array[8556]=30'd794287561;
array[8557]=30'd842495488;
array[8558]=30'd884420162;
array[8559]=30'd900139626;
array[8560]=30'd900139626;
array[8561]=30'd900139626;
array[8562]=30'd900139626;
array[8563]=30'd900139626;
array[8564]=30'd900139626;
array[8565]=30'd900139626;
array[8566]=30'd900139626;
array[8567]=30'd900139626;
array[8568]=30'd900139626;
array[8569]=30'd900139626;
array[8570]=30'd900139626;
array[8571]=30'd900139626;
array[8572]=30'd900139626;
array[8573]=30'd900139626;
array[8574]=30'd920102487;
array[8575]=30'd851962439;
array[8576]=30'd819475993;
array[8577]=30'd819475993;
array[8578]=30'd832058842;
array[8579]=30'd832058842;
array[8580]=30'd832058842;
array[8581]=30'd855119352;
array[8582]=30'd946320871;
array[8583]=30'd916923947;
array[8584]=30'd900139626;
array[8585]=30'd900139626;
array[8586]=30'd683036269;
array[8587]=30'd634745492;
array[8588]=30'd608524977;
array[8589]=30'd452327079;
array[8590]=30'd368466587;
array[8591]=30'd306613855;
array[8592]=30'd374749802;
array[8593]=30'd447089265;
array[8594]=30'd409379461;
array[8595]=30'd258398808;
array[8596]=30'd447089265;
array[8597]=30'd447089265;
array[8598]=30'd433483392;
array[8599]=30'd397823583;
array[8600]=30'd274187850;
array[8601]=30'd355962430;
array[8602]=30'd756500033;
array[8603]=30'd820432476;
array[8604]=30'd820432476;
array[8605]=30'd820432476;
array[8606]=30'd710361687;
array[8607]=30'd453521981;
array[8608]=30'd274187850;
array[8609]=30'd300461633;
array[8610]=30'd300461633;
array[8611]=30'd300461633;
array[8612]=30'd335980112;
array[8613]=30'd447089265;
array[8614]=30'd548772504;
array[8615]=30'd427157133;
array[8616]=30'd260455061;
array[8617]=30'd397823583;
array[8618]=30'd351684214;
array[8619]=30'd397823583;
array[8620]=30'd496374434;
array[8621]=30'd548772504;
array[8622]=30'd734429821;
array[8623]=30'd900139626;
array[8624]=30'd900139626;
array[8625]=30'd900139626;
array[8626]=30'd900139626;
array[8627]=30'd920102487;
array[8628]=30'd875032088;
array[8629]=30'd819475993;
array[8630]=30'd819437027;
array[8631]=30'd819437027;
array[8632]=30'd842495488;
array[8633]=30'd860306981;
array[8634]=30'd884420162;
array[8635]=30'd900139626;
array[8636]=30'd873911932;
array[8637]=30'd873911932;
array[8638]=30'd873911932;
array[8639]=30'd873911932;
array[8640]=30'd900139626;
array[8641]=30'd900139626;
array[8642]=30'd900139626;
array[8643]=30'd900139626;
array[8644]=30'd900139626;
array[8645]=30'd920102487;
array[8646]=30'd963075636;
array[8647]=30'd915924476;
array[8648]=30'd855119352;
array[8649]=30'd875032088;
array[8650]=30'd936883742;
array[8651]=30'd1016593896;
array[8652]=30'd926409165;
array[8653]=30'd794287561;
array[8654]=30'd884422147;
array[8655]=30'd916923947;
array[8656]=30'd900139626;
array[8657]=30'd898096696;
array[8658]=30'd851962439;
array[8659]=30'd851962439;
array[8660]=30'd884420162;
array[8661]=30'd900139626;
array[8662]=30'd900139626;
array[8663]=30'd900139626;
array[8664]=30'd900139626;
array[8665]=30'd900139626;
array[8666]=30'd900139626;
array[8667]=30'd900139626;
array[8668]=30'd900139626;
array[8669]=30'd920102487;
array[8670]=30'd851962439;
array[8671]=30'd819475993;
array[8672]=30'd983039487;
array[8673]=30'd963129822;
array[8674]=30'd963129822;
array[8675]=30'd946320871;
array[8676]=30'd896012764;
array[8677]=30'd819437027;
array[8678]=30'd915924476;
array[8679]=30'd916923947;
array[8680]=30'd900139626;
array[8681]=30'd900139626;
array[8682]=30'd625394265;
array[8683]=30'd634745492;
array[8684]=30'd591795877;
array[8685]=30'd427157133;
array[8686]=30'd351684214;
array[8687]=30'd335980112;
array[8688]=30'd351684214;
array[8689]=30'd447089265;
array[8690]=30'd409379461;
array[8691]=30'd258398808;
array[8692]=30'd447089265;
array[8693]=30'd456562280;
array[8694]=30'd385288799;
array[8695]=30'd294099551;
array[8696]=30'd300461633;
array[8697]=30'd409485846;
array[8698]=30'd710361687;
array[8699]=30'd820432476;
array[8700]=30'd803707487;
array[8701]=30'd589750888;
array[8702]=30'd274187850;
array[8703]=30'd300461633;
array[8704]=30'd282664514;
array[8705]=30'd282664514;
array[8706]=30'd300461633;
array[8707]=30'd300461633;
array[8708]=30'd335980112;
array[8709]=30'd559296136;
array[8710]=30'd461756049;
array[8711]=30'd368466587;
array[8712]=30'd277255789;
array[8713]=30'd456562280;
array[8714]=30'd306613855;
array[8715]=30'd397823583;
array[8716]=30'd461756049;
array[8717]=30'd525726362;
array[8718]=30'd791076458;
array[8719]=30'd900139626;
array[8720]=30'd900139626;
array[8721]=30'd900139626;
array[8722]=30'd900139626;
array[8723]=30'd900139626;
array[8724]=30'd900139626;
array[8725]=30'd900139626;
array[8726]=30'd884420162;
array[8727]=30'd884420162;
array[8728]=30'd884420162;
array[8729]=30'd884420162;
array[8730]=30'd900139626;
array[8731]=30'd900139626;
array[8732]=30'd873911932;
array[8733]=30'd873911932;
array[8734]=30'd873911932;
array[8735]=30'd873911932;
array[8736]=30'd900139626;
array[8737]=30'd900139626;
array[8738]=30'd900139626;
array[8739]=30'd900139626;
array[8740]=30'd900139626;
array[8741]=30'd920102487;
array[8742]=30'd875032088;
array[8743]=30'd785935846;
array[8744]=30'd785935846;
array[8745]=30'd785935846;
array[8746]=30'd785935846;
array[8747]=30'd946320871;
array[8748]=30'd983039487;
array[8749]=30'd896012764;
array[8750]=30'd819437027;
array[8751]=30'd884422147;
array[8752]=30'd898096696;
array[8753]=30'd819475993;
array[8754]=30'd785935846;
array[8755]=30'd842495488;
array[8756]=30'd884420162;
array[8757]=30'd900139626;
array[8758]=30'd900139626;
array[8759]=30'd900139626;
array[8760]=30'd900139626;
array[8761]=30'd900139626;
array[8762]=30'd900139626;
array[8763]=30'd900139626;
array[8764]=30'd920102487;
array[8765]=30'd851962439;
array[8766]=30'd855119352;
array[8767]=30'd963129822;
array[8768]=30'd963129822;
array[8769]=30'd896012764;
array[8770]=30'd855119352;
array[8771]=30'd832058842;
array[8772]=30'd870853059;
array[8773]=30'd832058842;
array[8774]=30'd832058842;
array[8775]=30'd916923947;
array[8776]=30'd900139626;
array[8777]=30'd900139626;
array[8778]=30'd625394265;
array[8779]=30'd634745492;
array[8780]=30'd591795877;
array[8781]=30'd409379461;
array[8782]=30'd351684214;
array[8783]=30'd374749802;
array[8784]=30'd333912689;
array[8785]=30'd447089265;
array[8786]=30'd456562280;
array[8787]=30'd335980112;
array[8788]=30'd363288160;
array[8789]=30'd312961612;
array[8790]=30'd274187850;
array[8791]=30'd300461633;
array[8792]=30'd300461633;
array[8793]=30'd407406158;
array[8794]=30'd778553911;
array[8795]=30'd778553911;
array[8796]=30'd453521981;
array[8797]=30'd274187850;
array[8798]=30'd300461633;
array[8799]=30'd282664514;
array[8800]=30'd282664514;
array[8801]=30'd282664514;
array[8802]=30'd300461633;
array[8803]=30'd234392123;
array[8804]=30'd456562280;
array[8805]=30'd525726362;
array[8806]=30'd427157133;
array[8807]=30'd306613855;
array[8808]=30'd385288799;
array[8809]=30'd456562280;
array[8810]=30'd306613855;
array[8811]=30'd397823583;
array[8812]=30'd461756049;
array[8813]=30'd525726362;
array[8814]=30'd791076458;
array[8815]=30'd900139626;
array[8816]=30'd900139626;
array[8817]=30'd900139626;
array[8818]=30'd900139626;
array[8819]=30'd900139626;
array[8820]=30'd900139626;
array[8821]=30'd900139626;
array[8822]=30'd900139626;
array[8823]=30'd900139626;
array[8824]=30'd900139626;
array[8825]=30'd900139626;
array[8826]=30'd900139626;
array[8827]=30'd900139626;
array[8828]=30'd873911932;
array[8829]=30'd873911932;
array[8830]=30'd873911932;
array[8831]=30'd873911932;
array[8832]=30'd900139626;
array[8833]=30'd900139626;
array[8834]=30'd900139626;
array[8835]=30'd900139626;
array[8836]=30'd900139626;
array[8837]=30'd920102487;
array[8838]=30'd819475993;
array[8839]=30'd894973365;
array[8840]=30'd944268729;
array[8841]=30'd914919842;
array[8842]=30'd778588583;
array[8843]=30'd832058842;
array[8844]=30'd946320871;
array[8845]=30'd963129822;
array[8846]=30'd794287561;
array[8847]=30'd884422147;
array[8848]=30'd936883742;
array[8849]=30'd983039487;
array[8850]=30'd983039487;
array[8851]=30'd916923947;
array[8852]=30'd884420162;
array[8853]=30'd900139626;
array[8854]=30'd900139626;
array[8855]=30'd900139626;
array[8856]=30'd900139626;
array[8857]=30'd900139626;
array[8858]=30'd900139626;
array[8859]=30'd900139626;
array[8860]=30'd898096696;
array[8861]=30'd819475993;
array[8862]=30'd963129822;
array[8863]=30'd963129822;
array[8864]=30'd776468978;
array[8865]=30'd670582270;
array[8866]=30'd670582270;
array[8867]=30'd650619404;
array[8868]=30'd635956692;
array[8869]=30'd541577678;
array[8870]=30'd754446794;
array[8871]=30'd963077644;
array[8872]=30'd884420162;
array[8873]=30'd900139626;
array[8874]=30'd589750888;
array[8875]=30'd634745492;
array[8876]=30'd548772504;
array[8877]=30'd328601227;
array[8878]=30'd306613855;
array[8879]=30'd421932631;
array[8880]=30'd363288160;
array[8881]=30'd333912689;
array[8882]=30'd363288160;
array[8883]=30'd274187850;
array[8884]=30'd247985748;
array[8885]=30'd234392123;
array[8886]=30'd300461633;
array[8887]=30'd300461633;
array[8888]=30'd282664514;
array[8889]=30'd340285012;
array[8890]=30'd726149706;
array[8891]=30'd407406158;
array[8892]=30'd234392123;
array[8893]=30'd300461633;
array[8894]=30'd282664514;
array[8895]=30'd282664514;
array[8896]=30'd282664514;
array[8897]=30'd282664514;
array[8898]=30'd300461633;
array[8899]=30'd274187850;
array[8900]=30'd559296136;
array[8901]=30'd461756049;
array[8902]=30'd368466587;
array[8903]=30'd234283624;
array[8904]=30'd277255789;
array[8905]=30'd363288160;
array[8906]=30'd306613855;
array[8907]=30'd374749802;
array[8908]=30'd484819572;
array[8909]=30'd525726362;
array[8910]=30'd820432476;
array[8911]=30'd900139626;
array[8912]=30'd900139626;
array[8913]=30'd900139626;
array[8914]=30'd900139626;
array[8915]=30'd900139626;
array[8916]=30'd900139626;
array[8917]=30'd900139626;
array[8918]=30'd900139626;
array[8919]=30'd900139626;
array[8920]=30'd900139626;
array[8921]=30'd900139626;
array[8922]=30'd900139626;
array[8923]=30'd900139626;
array[8924]=30'd900139626;
array[8925]=30'd900139626;
array[8926]=30'd900139626;
array[8927]=30'd900139626;
array[8928]=30'd900139626;
array[8929]=30'd900139626;
array[8930]=30'd900139626;
array[8931]=30'd900139626;
array[8932]=30'd920102487;
array[8933]=30'd898096696;
array[8934]=30'd785935846;
array[8935]=30'd894973365;
array[8936]=30'd854099361;
array[8937]=30'd914919842;
array[8938]=30'd870853059;
array[8939]=30'd810051001;
array[8940]=30'd915924476;
array[8941]=30'd963129822;
array[8942]=30'd794287561;
array[8943]=30'd884422147;
array[8944]=30'd915924476;
array[8945]=30'd915924476;
array[8946]=30'd915924476;
array[8947]=30'd916923947;
array[8948]=30'd916923947;
array[8949]=30'd900139626;
array[8950]=30'd900139626;
array[8951]=30'd900139626;
array[8952]=30'd900139626;
array[8953]=30'd900139626;
array[8954]=30'd900139626;
array[8955]=30'd900139626;
array[8956]=30'd898096696;
array[8957]=30'd819475993;
array[8958]=30'd855119352;
array[8959]=30'd708318695;
array[8960]=30'd708318695;
array[8961]=30'd896012764;
array[8962]=30'd963129822;
array[8963]=30'd983039487;
array[8964]=30'd946320871;
array[8965]=30'd708318695;
array[8966]=30'd690495950;
array[8967]=30'd946320871;
array[8968]=30'd884420162;
array[8969]=30'd900139626;
array[8970]=30'd556154453;
array[8971]=30'd634745492;
array[8972]=30'd525726362;
array[8973]=30'd300284569;
array[8974]=30'd277255789;
array[8975]=30'd363288160;
array[8976]=30'd407406158;
array[8977]=30'd453540449;
array[8978]=30'd453540449;
array[8979]=30'd315184704;
array[8980]=30'd282664514;
array[8981]=30'd239672891;
array[8982]=30'd282664514;
array[8983]=30'd282664514;
array[8984]=30'd282664514;
array[8985]=30'd254351946;
array[8986]=30'd340285012;
array[8987]=30'd279466521;
array[8988]=30'd300461633;
array[8989]=30'd282664514;
array[8990]=30'd282664514;
array[8991]=30'd282664514;
array[8992]=30'd282664514;
array[8993]=30'd282664514;
array[8994]=30'd234392123;
array[8995]=30'd484874837;
array[8996]=30'd503733877;
array[8997]=30'd433483392;
array[8998]=30'd260455061;
array[8999]=30'd234283624;
array[9000]=30'd274187850;
array[9001]=30'd247985748;
array[9002]=30'd220707388;
array[9003]=30'd335980112;
array[9004]=30'd447089265;
array[9005]=30'd503733877;
array[9006]=30'd791076458;
array[9007]=30'd900139626;
array[9008]=30'd873911932;
array[9009]=30'd900139626;
array[9010]=30'd900139626;
array[9011]=30'd900139626;
array[9012]=30'd900139626;
array[9013]=30'd900139626;
array[9014]=30'd900139626;
array[9015]=30'd900139626;
array[9016]=30'd900139626;
array[9017]=30'd900139626;
array[9018]=30'd900139626;
array[9019]=30'd900139626;
array[9020]=30'd900139626;
array[9021]=30'd900139626;
array[9022]=30'd900139626;
array[9023]=30'd900139626;
array[9024]=30'd860306981;
array[9025]=30'd884420162;
array[9026]=30'd900139626;
array[9027]=30'd900139626;
array[9028]=30'd920102487;
array[9029]=30'd875032088;
array[9030]=30'd810051001;
array[9031]=30'd854099361;
array[9032]=30'd790145435;
array[9033]=30'd914919842;
array[9034]=30'd914919842;
array[9035]=30'd810051001;
array[9036]=30'd896012764;
array[9037]=30'd963129822;
array[9038]=30'd794287561;
array[9039]=30'd896012764;
array[9040]=30'd855119352;
array[9041]=30'd785935846;
array[9042]=30'd785935846;
array[9043]=30'd842495488;
array[9044]=30'd916923947;
array[9045]=30'd900139626;
array[9046]=30'd900139626;
array[9047]=30'd900139626;
array[9048]=30'd900139626;
array[9049]=30'd900139626;
array[9050]=30'd900139626;
array[9051]=30'd851962439;
array[9052]=30'd728246811;
array[9053]=30'd751308299;
array[9054]=30'd915924476;
array[9055]=30'd1034407430;
array[9056]=30'd1034407430;
array[9057]=30'd1034407430;
array[9058]=30'd1034407430;
array[9059]=30'd1034407430;
array[9060]=30'd1016593896;
array[9061]=30'd875032088;
array[9062]=30'd581437943;
array[9063]=30'd963077644;
array[9064]=30'd941029952;
array[9065]=30'd900139626;
array[9066]=30'd530993763;
array[9067]=30'd634745492;
array[9068]=30'd525726362;
array[9069]=30'd260455061;
array[9070]=30'd340285012;
array[9071]=30'd481853012;
array[9072]=30'd473528913;
array[9073]=30'd473528913;
array[9074]=30'd473528913;
array[9075]=30'd414803529;
array[9076]=30'd282664514;
array[9077]=30'd239672891;
array[9078]=30'd282664514;
array[9079]=30'd282664514;
array[9080]=30'd282664514;
array[9081]=30'd239672891;
array[9082]=30'd254351946;
array[9083]=30'd300461633;
array[9084]=30'd282664514;
array[9085]=30'd282664514;
array[9086]=30'd282664514;
array[9087]=30'd282664514;
array[9088]=30'd282664514;
array[9089]=30'd300461633;
array[9090]=30'd312961612;
array[9091]=30'd556154453;
array[9092]=30'd427157133;
array[9093]=30'd368466587;
array[9094]=30'd294099551;
array[9095]=30'd274187850;
array[9096]=30'd340285012;
array[9097]=30'd352935499;
array[9098]=30'd381210191;
array[9099]=30'd340285012;
array[9100]=30'd363288160;
array[9101]=30'd503733877;
array[9102]=30'd734429821;
array[9103]=30'd900139626;
array[9104]=30'd900139626;
array[9105]=30'd900139626;
array[9106]=30'd900139626;
array[9107]=30'd900139626;
array[9108]=30'd900139626;
array[9109]=30'd900139626;
array[9110]=30'd900139626;
array[9111]=30'd900139626;
array[9112]=30'd900139626;
array[9113]=30'd900139626;
array[9114]=30'd900139626;
array[9115]=30'd900139626;
array[9116]=30'd900139626;
array[9117]=30'd900139626;
array[9118]=30'd900139626;
array[9119]=30'd900139626;
array[9120]=30'd650619404;
array[9121]=30'd884420162;
array[9122]=30'd920102487;
array[9123]=30'd920102487;
array[9124]=30'd920102487;
array[9125]=30'd875032088;
array[9126]=30'd810051001;
array[9127]=30'd883468684;
array[9128]=30'd810051001;
array[9129]=30'd914919842;
array[9130]=30'd914919842;
array[9131]=30'd764966339;
array[9132]=30'd896012764;
array[9133]=30'd896012764;
array[9134]=30'd794287561;
array[9135]=30'd946320871;
array[9136]=30'd946320871;
array[9137]=30'd915924476;
array[9138]=30'd896012764;
array[9139]=30'd842495488;
array[9140]=30'd916923947;
array[9141]=30'd916923947;
array[9142]=30'd884420162;
array[9143]=30'd884420162;
array[9144]=30'd884420162;
array[9145]=30'd839339599;
array[9146]=30'd710361687;
array[9147]=30'd778553911;
array[9148]=30'd936883742;
array[9149]=30'd1034407430;
array[9150]=30'd1034407430;
array[9151]=30'd1034407430;
array[9152]=30'd1034407430;
array[9153]=30'd1034407430;
array[9154]=30'd1034407430;
array[9155]=30'd1034407430;
array[9156]=30'd1034407430;
array[9157]=30'd842495488;
array[9158]=30'd503787028;
array[9159]=30'd793183798;
array[9160]=30'd900139626;
array[9161]=30'd900139626;
array[9162]=30'd568785526;
array[9163]=30'd634745492;
array[9164]=30'd496374434;
array[9165]=30'd277255789;
array[9166]=30'd432564808;
array[9167]=30'd518575683;
array[9168]=30'd473528913;
array[9169]=30'd473528913;
array[9170]=30'd473528913;
array[9171]=30'd458840642;
array[9172]=30'd315184704;
array[9173]=30'd254351946;
array[9174]=30'd282664514;
array[9175]=30'd282664514;
array[9176]=30'd282664514;
array[9177]=30'd239672891;
array[9178]=30'd206118464;
array[9179]=30'd282664514;
array[9180]=30'd282664514;
array[9181]=30'd282664514;
array[9182]=30'd282664514;
array[9183]=30'd282664514;
array[9184]=30'd282664514;
array[9185]=30'd300461633;
array[9186]=30'd456562280;
array[9187]=30'd503733877;
array[9188]=30'd427157133;
array[9189]=30'd333912689;
array[9190]=30'd363288160;
array[9191]=30'd432564808;
array[9192]=30'd458840642;
array[9193]=30'd458840642;
array[9194]=30'd458840642;
array[9195]=30'd494467625;
array[9196]=30'd432564808;
array[9197]=30'd421987917;
array[9198]=30'd710361687;
array[9199]=30'd900139626;
array[9200]=30'd900139626;
array[9201]=30'd900139626;
array[9202]=30'd900139626;
array[9203]=30'd900139626;
array[9204]=30'd900139626;
array[9205]=30'd900139626;
array[9206]=30'd900139626;
array[9207]=30'd900139626;
array[9208]=30'd900139626;
array[9209]=30'd900139626;
array[9210]=30'd900139626;
array[9211]=30'd900139626;
array[9212]=30'd900139626;
array[9213]=30'd900139626;
array[9214]=30'd900139626;
array[9215]=30'd900139626;
array[9216]=30'd465022394;
array[9217]=30'd724009508;
array[9218]=30'd920102487;
array[9219]=30'd920102487;
array[9220]=30'd920102487;
array[9221]=30'd915924476;
array[9222]=30'd810051001;
array[9223]=30'd854099361;
array[9224]=30'd790145435;
array[9225]=30'd790145435;
array[9226]=30'd810051001;
array[9227]=30'd870853059;
array[9228]=30'd926409165;
array[9229]=30'd870853059;
array[9230]=30'd832058842;
array[9231]=30'd896012764;
array[9232]=30'd946320871;
array[9233]=30'd983039487;
array[9234]=30'd963077644;
array[9235]=30'd936883742;
array[9236]=30'd884420162;
array[9237]=30'd756500033;
array[9238]=30'd756500033;
array[9239]=30'd860306981;
array[9240]=30'd860306981;
array[9241]=30'd681011766;
array[9242]=30'd681011766;
array[9243]=30'd936883742;
array[9244]=30'd1002945052;
array[9245]=30'd1034407430;
array[9246]=30'd1034407430;
array[9247]=30'd1034407430;
array[9248]=30'd1034407430;
array[9249]=30'd1002945052;
array[9250]=30'd1034407430;
array[9251]=30'd1002945052;
array[9252]=30'd936883742;
array[9253]=30'd556235306;
array[9254]=30'd756500033;
array[9255]=30'd941029952;
array[9256]=30'd900139626;
array[9257]=30'd900139626;
array[9258]=30'd589750888;
array[9259]=30'd650530435;
array[9260]=30'd474371718;
array[9261]=30'd294099551;
array[9262]=30'd453540449;
array[9263]=30'd473528913;
array[9264]=30'd473528913;
array[9265]=30'd473528913;
array[9266]=30'd473528913;
array[9267]=30'd473528913;
array[9268]=30'd352935499;
array[9269]=30'd282664514;
array[9270]=30'd282664514;
array[9271]=30'd282664514;
array[9272]=30'd239672891;
array[9273]=30'd239672891;
array[9274]=30'd206118464;
array[9275]=30'd239672891;
array[9276]=30'd282664514;
array[9277]=30'd282664514;
array[9278]=30'd282664514;
array[9279]=30'd282664514;
array[9280]=30'd282664514;
array[9281]=30'd274187850;
array[9282]=30'd530993763;
array[9283]=30'd433483392;
array[9284]=30'd368466587;
array[9285]=30'd385288799;
array[9286]=30'd363288160;
array[9287]=30'd481853012;
array[9288]=30'd458840642;
array[9289]=30'd473528913;
array[9290]=30'd473528913;
array[9291]=30'd473528913;
array[9292]=30'd458840642;
array[9293]=30'd432564808;
array[9294]=30'd586701367;
array[9295]=30'd920102487;
array[9296]=30'd900139626;
array[9297]=30'd900139626;
array[9298]=30'd900139626;
array[9299]=30'd900139626;
array[9300]=30'd900139626;
array[9301]=30'd900139626;
array[9302]=30'd900139626;
array[9303]=30'd900139626;
array[9304]=30'd900139626;
array[9305]=30'd900139626;
array[9306]=30'd900139626;
array[9307]=30'd900139626;
array[9308]=30'd900139626;
array[9309]=30'd900139626;
array[9310]=30'd900139626;
array[9311]=30'd900139626;
array[9312]=30'd478665137;
array[9313]=30'd489151968;
array[9314]=30'd808945195;
array[9315]=30'd920102487;
array[9316]=30'd920102487;
array[9317]=30'd963075636;
array[9318]=30'd896012764;
array[9319]=30'd790145435;
array[9320]=30'd854099361;
array[9321]=30'd883468684;
array[9322]=30'd914919842;
array[9323]=30'd894973365;
array[9324]=30'd810051001;
array[9325]=30'd810051001;
array[9326]=30'd832058842;
array[9327]=30'd776468978;
array[9328]=30'd819437027;
array[9329]=30'd842495488;
array[9330]=30'd860306981;
array[9331]=30'd778553911;
array[9332]=30'd724009508;
array[9333]=30'd884420162;
array[9334]=30'd963075636;
array[9335]=30'd963075636;
array[9336]=30'd963075636;
array[9337]=30'd963075636;
array[9338]=30'd778553911;
array[9339]=30'd724009508;
array[9340]=30'd936883742;
array[9341]=30'd1002945052;
array[9342]=30'd963077644;
array[9343]=30'd875032088;
array[9344]=30'd808945195;
array[9345]=30'd751308299;
array[9346]=30'd778553911;
array[9347]=30'd756500033;
array[9348]=30'd808945195;
array[9349]=30'd839339599;
array[9350]=30'd574048834;
array[9351]=30'd839339599;
array[9352]=30'd900139626;
array[9353]=30'd900139626;
array[9354]=30'd547846737;
array[9355]=30'd625322602;
array[9356]=30'd503733877;
array[9357]=30'd294099551;
array[9358]=30'd481853012;
array[9359]=30'd473528913;
array[9360]=30'd488205898;
array[9361]=30'd488205898;
array[9362]=30'd473528913;
array[9363]=30'd473528913;
array[9364]=30'd414803529;
array[9365]=30'd282664514;
array[9366]=30'd254351946;
array[9367]=30'd239672891;
array[9368]=30'd206118464;
array[9369]=30'd206118464;
array[9370]=30'd239672891;
array[9371]=30'd239672891;
array[9372]=30'd254351946;
array[9373]=30'd282664514;
array[9374]=30'd315184704;
array[9375]=30'd315184704;
array[9376]=30'd415828509;
array[9377]=30'd355962430;
array[9378]=30'd559296136;
array[9379]=30'd433483392;
array[9380]=30'd277255789;
array[9381]=30'd421987917;
array[9382]=30'd340285012;
array[9383]=30'd481853012;
array[9384]=30'd473528913;
array[9385]=30'd473528913;
array[9386]=30'd473528913;
array[9387]=30'd473528913;
array[9388]=30'd414803529;
array[9389]=30'd414803529;
array[9390]=30'd432564808;
array[9391]=30'd803707487;
array[9392]=30'd900139626;
array[9393]=30'd900139626;
array[9394]=30'd900139626;
array[9395]=30'd900139626;
array[9396]=30'd900139626;
array[9397]=30'd900139626;
array[9398]=30'd900139626;
array[9399]=30'd900139626;
array[9400]=30'd900139626;
array[9401]=30'd900139626;
array[9402]=30'd900139626;
array[9403]=30'd900139626;
array[9404]=30'd900139626;
array[9405]=30'd900139626;
array[9406]=30'd900139626;
array[9407]=30'd900139626;
array[9408]=30'd478665137;
array[9409]=30'd465022394;
array[9410]=30'd520605190;
array[9411]=30'd851962439;
array[9412]=30'd920102487;
array[9413]=30'd963075636;
array[9414]=30'd983039487;
array[9415]=30'd810051001;
array[9416]=30'd790145435;
array[9417]=30'd854099361;
array[9418]=30'd790145435;
array[9419]=30'd810051001;
array[9420]=30'd870853059;
array[9421]=30'd896012764;
array[9422]=30'd963129822;
array[9423]=30'd776468978;
array[9424]=30'd691505656;
array[9425]=30'd808945195;
array[9426]=30'd613919272;
array[9427]=30'd808945195;
array[9428]=30'd963075636;
array[9429]=30'd963075636;
array[9430]=30'd963075636;
array[9431]=30'd963075636;
array[9432]=30'd963075636;
array[9433]=30'd963075636;
array[9434]=30'd963075636;
array[9435]=30'd613919272;
array[9436]=30'd598167087;
array[9437]=30'd724009508;
array[9438]=30'd808945195;
array[9439]=30'd860306981;
array[9440]=30'd898096696;
array[9441]=30'd920102487;
array[9442]=30'd898096696;
array[9443]=30'd920102487;
array[9444]=30'd941029952;
array[9445]=30'd920102487;
array[9446]=30'd900139626;
array[9447]=30'd900139626;
array[9448]=30'd900139626;
array[9449]=30'd803707487;
array[9450]=30'd363288160;
array[9451]=30'd556154453;
array[9452]=30'd503733877;
array[9453]=30'd294099551;
array[9454]=30'd518575683;
array[9455]=30'd473528913;
array[9456]=30'd473528913;
array[9457]=30'd488205898;
array[9458]=30'd473528913;
array[9459]=30'd473528913;
array[9460]=30'd458840642;
array[9461]=30'd315184704;
array[9462]=30'd315184704;
array[9463]=30'd282664514;
array[9464]=30'd239672891;
array[9465]=30'd206118464;
array[9466]=30'd282664514;
array[9467]=30'd315184704;
array[9468]=30'd282664514;
array[9469]=30'd352935499;
array[9470]=30'd458840642;
array[9471]=30'd414803529;
array[9472]=30'd371776054;
array[9473]=30'd421987917;
array[9474]=30'd503733877;
array[9475]=30'd385288799;
array[9476]=30'd199687791;
array[9477]=30'd363288160;
array[9478]=30'd407406158;
array[9479]=30'd481853012;
array[9480]=30'd473528913;
array[9481]=30'd473528913;
array[9482]=30'd473528913;
array[9483]=30'd458840642;
array[9484]=30'd414803529;
array[9485]=30'd473528913;
array[9486]=30'd458840642;
array[9487]=30'd565736011;
array[9488]=30'd920102487;
array[9489]=30'd900139626;
array[9490]=30'd900139626;
array[9491]=30'd900139626;
array[9492]=30'd900139626;
array[9493]=30'd900139626;
array[9494]=30'd900139626;
array[9495]=30'd900139626;
array[9496]=30'd900139626;
array[9497]=30'd900139626;
array[9498]=30'd900139626;
array[9499]=30'd900139626;
array[9500]=30'd900139626;
array[9501]=30'd900139626;
array[9502]=30'd900139626;
array[9503]=30'd900139626;
array[9504]=30'd478665137;
array[9505]=30'd465022394;
array[9506]=30'd465022394;
array[9507]=30'd650619404;
array[9508]=30'd898096696;
array[9509]=30'd920102487;
array[9510]=30'd1002945052;
array[9511]=30'd963129822;
array[9512]=30'd870853059;
array[9513]=30'd870853059;
array[9514]=30'd926409165;
array[9515]=30'd946320871;
array[9516]=30'd915924476;
array[9517]=30'd936883742;
array[9518]=30'd778553911;
array[9519]=30'd860306981;
array[9520]=30'd936883742;
array[9521]=30'd963077644;
array[9522]=30'd724009508;
array[9523]=30'd916923947;
array[9524]=30'd963075636;
array[9525]=30'd963075636;
array[9526]=30'd963075636;
array[9527]=30'd963075636;
array[9528]=30'd963075636;
array[9529]=30'd963075636;
array[9530]=30'd963075636;
array[9531]=30'd808945195;
array[9532]=30'd839339599;
array[9533]=30'd920102487;
array[9534]=30'd920102487;
array[9535]=30'd920102487;
array[9536]=30'd920102487;
array[9537]=30'd920102487;
array[9538]=30'd920102487;
array[9539]=30'd920102487;
array[9540]=30'd900139626;
array[9541]=30'd900139626;
array[9542]=30'd900139626;
array[9543]=30'd920102487;
array[9544]=30'd900139626;
array[9545]=30'd565736011;
array[9546]=30'd453521981;
array[9547]=30'd456562280;
array[9548]=30'd503733877;
array[9549]=30'd355962430;
array[9550]=30'd518575683;
array[9551]=30'd473528913;
array[9552]=30'd488205898;
array[9553]=30'd488205898;
array[9554]=30'd488205898;
array[9555]=30'd473528913;
array[9556]=30'd488205898;
array[9557]=30'd473528913;
array[9558]=30'd458840642;
array[9559]=30'd458840642;
array[9560]=30'd415828509;
array[9561]=30'd282664514;
array[9562]=30'd414803529;
array[9563]=30'd458840642;
array[9564]=30'd458840642;
array[9565]=30'd414803529;
array[9566]=30'd414803529;
array[9567]=30'd352935499;
array[9568]=30'd432564808;
array[9569]=30'd470243883;
array[9570]=30'd456562280;
array[9571]=30'd294099551;
array[9572]=30'd224918107;
array[9573]=30'd340285012;
array[9574]=30'd432564808;
array[9575]=30'd481853012;
array[9576]=30'd473528913;
array[9577]=30'd473528913;
array[9578]=30'd458840642;
array[9579]=30'd414803529;
array[9580]=30'd458840642;
array[9581]=30'd473528913;
array[9582]=30'd473528913;
array[9583]=30'd414803529;
array[9584]=30'd851962439;
array[9585]=30'd920102487;
array[9586]=30'd900139626;
array[9587]=30'd900139626;
array[9588]=30'd900139626;
array[9589]=30'd900139626;
array[9590]=30'd900139626;
array[9591]=30'd900139626;
array[9592]=30'd900139626;
array[9593]=30'd900139626;
array[9594]=30'd900139626;
array[9595]=30'd900139626;
array[9596]=30'd900139626;
array[9597]=30'd900139626;
array[9598]=30'd900139626;
array[9599]=30'd900139626;
array[9600]=30'd445105582;
array[9601]=30'd465022394;
array[9602]=30'd445105582;
array[9603]=30'd405258689;
array[9604]=30'd650619404;
array[9605]=30'd728246811;
array[9606]=30'd778553911;
array[9607]=30'd819475993;
array[9608]=30'd776468978;
array[9609]=30'd776468978;
array[9610]=30'd875032088;
array[9611]=30'd936883742;
array[9612]=30'd898096696;
array[9613]=30'd920102487;
array[9614]=30'd756500033;
array[9615]=30'd936883742;
array[9616]=30'd936883742;
array[9617]=30'd778553911;
array[9618]=30'd860306981;
array[9619]=30'd963075636;
array[9620]=30'd963075636;
array[9621]=30'd963075636;
array[9622]=30'd963075636;
array[9623]=30'd963075636;
array[9624]=30'd963075636;
array[9625]=30'd963075636;
array[9626]=30'd963075636;
array[9627]=30'd884420162;
array[9628]=30'd839339599;
array[9629]=30'd920102487;
array[9630]=30'd920102487;
array[9631]=30'd920102487;
array[9632]=30'd920102487;
array[9633]=30'd920102487;
array[9634]=30'd920102487;
array[9635]=30'd920102487;
array[9636]=30'd920102487;
array[9637]=30'd900139626;
array[9638]=30'd920102487;
array[9639]=30'd920102487;
array[9640]=30'd782746219;
array[9641]=30'd453540449;
array[9642]=30'd481853012;
array[9643]=30'd407406158;
array[9644]=30'd506984008;
array[9645]=30'd340285012;
array[9646]=30'd481853012;
array[9647]=30'd473528913;
array[9648]=30'd488205898;
array[9649]=30'd488205898;
array[9650]=30'd488205898;
array[9651]=30'd488205898;
array[9652]=30'd488205898;
array[9653]=30'd473528913;
array[9654]=30'd473528913;
array[9655]=30'd473528913;
array[9656]=30'd458840642;
array[9657]=30'd414803529;
array[9658]=30'd473528913;
array[9659]=30'd473528913;
array[9660]=30'd473528913;
array[9661]=30'd473528913;
array[9662]=30'd473528913;
array[9663]=30'd458840642;
array[9664]=30'd458840642;
array[9665]=30'd421987917;
array[9666]=30'd456562280;
array[9667]=30'd294099551;
array[9668]=30'd407406158;
array[9669]=30'd300461633;
array[9670]=30'd432564808;
array[9671]=30'd473528913;
array[9672]=30'd473528913;
array[9673]=30'd473528913;
array[9674]=30'd414803529;
array[9675]=30'd458840642;
array[9676]=30'd473528913;
array[9677]=30'd473528913;
array[9678]=30'd473528913;
array[9679]=30'd458840642;
array[9680]=30'd698886706;
array[9681]=30'd920102487;
array[9682]=30'd900139626;
array[9683]=30'd900139626;
array[9684]=30'd900139626;
array[9685]=30'd900139626;
array[9686]=30'd900139626;
array[9687]=30'd900139626;
array[9688]=30'd900139626;
array[9689]=30'd900139626;
array[9690]=30'd900139626;
array[9691]=30'd900139626;
array[9692]=30'd900139626;
array[9693]=30'd900139626;
array[9694]=30'd900139626;
array[9695]=30'd920102487;
array[9696]=30'd445105582;
array[9697]=30'd445105582;
array[9698]=30'd465022394;
array[9699]=30'd445105582;
array[9700]=30'd445105582;
array[9701]=30'd425177566;
array[9702]=30'd609741283;
array[9703]=30'd915924476;
array[9704]=30'd983039487;
array[9705]=30'd1002945052;
array[9706]=30'd920102487;
array[9707]=30'd920102487;
array[9708]=30'd920102487;
array[9709]=30'd920102487;
array[9710]=30'd803707487;
array[9711]=30'd641178184;
array[9712]=30'd756500033;
array[9713]=30'd936883742;
array[9714]=30'd963075636;
array[9715]=30'd963075636;
array[9716]=30'd963075636;
array[9717]=30'd963075636;
array[9718]=30'd963075636;
array[9719]=30'd963075636;
array[9720]=30'd963075636;
array[9721]=30'd963075636;
array[9722]=30'd963075636;
array[9723]=30'd860306981;
array[9724]=30'd839339599;
array[9725]=30'd920102487;
array[9726]=30'd920102487;
array[9727]=30'd920102487;
array[9728]=30'd920102487;
array[9729]=30'd920102487;
array[9730]=30'd920102487;
array[9731]=30'd920102487;
array[9732]=30'd920102487;
array[9733]=30'd920102487;
array[9734]=30'd920102487;
array[9735]=30'd851962439;
array[9736]=30'd506984008;
array[9737]=30'd518575683;
array[9738]=30'd473528913;
array[9739]=30'd481853012;
array[9740]=30'd340285012;
array[9741]=30'd340285012;
array[9742]=30'd381210191;
array[9743]=30'd458840642;
array[9744]=30'd488205898;
array[9745]=30'd488205898;
array[9746]=30'd488205898;
array[9747]=30'd488205898;
array[9748]=30'd488205898;
array[9749]=30'd473528913;
array[9750]=30'd473528913;
array[9751]=30'd473528913;
array[9752]=30'd414803529;
array[9753]=30'd473528913;
array[9754]=30'd473528913;
array[9755]=30'd488205898;
array[9756]=30'd488205898;
array[9757]=30'd473528913;
array[9758]=30'd473528913;
array[9759]=30'd473528913;
array[9760]=30'd458840642;
array[9761]=30'd340285012;
array[9762]=30'd340285012;
array[9763]=30'd407406158;
array[9764]=30'd481853012;
array[9765]=30'd371776054;
array[9766]=30'd381210191;
array[9767]=30'd473528913;
array[9768]=30'd473528913;
array[9769]=30'd458840642;
array[9770]=30'd414803529;
array[9771]=30'd473528913;
array[9772]=30'd473528913;
array[9773]=30'd473528913;
array[9774]=30'd473528913;
array[9775]=30'd458840642;
array[9776]=30'd565736011;
array[9777]=30'd920102487;
array[9778]=30'd900139626;
array[9779]=30'd900139626;
array[9780]=30'd900139626;
array[9781]=30'd900139626;
array[9782]=30'd900139626;
array[9783]=30'd900139626;
array[9784]=30'd920102487;
array[9785]=30'd920102487;
array[9786]=30'd920102487;
array[9787]=30'd920102487;
array[9788]=30'd920102487;
array[9789]=30'd920102487;
array[9790]=30'd920102487;
array[9791]=30'd920102487;
array[9792]=30'd465022394;
array[9793]=30'd465022394;
array[9794]=30'd478665137;
array[9795]=30'd465022394;
array[9796]=30'd478665137;
array[9797]=30'd491240873;
array[9798]=30'd776468978;
array[9799]=30'd983039487;
array[9800]=30'd983039487;
array[9801]=30'd1002945052;
array[9802]=30'd963075636;
array[9803]=30'd920102487;
array[9804]=30'd920102487;
array[9805]=30'd920102487;
array[9806]=30'd920102487;
array[9807]=30'd710361687;
array[9808]=30'd916923947;
array[9809]=30'd981941808;
array[9810]=30'd963075636;
array[9811]=30'd963075636;
array[9812]=30'd963075636;
array[9813]=30'd963075636;
array[9814]=30'd963075636;
array[9815]=30'd963075636;
array[9816]=30'd963075636;
array[9817]=30'd963075636;
array[9818]=30'd963075636;
array[9819]=30'd756500033;
array[9820]=30'd884420162;
array[9821]=30'd920102487;
array[9822]=30'd920102487;
array[9823]=30'd920102487;
array[9824]=30'd920102487;
array[9825]=30'd920102487;
array[9826]=30'd920102487;
array[9827]=30'd920102487;
array[9828]=30'd920102487;
array[9829]=30'd920102487;
array[9830]=30'd884420162;
array[9831]=30'd506984008;
array[9832]=30'd481853012;
array[9833]=30'd473528913;
array[9834]=30'd473528913;
array[9835]=30'd473528913;
array[9836]=30'd407406158;
array[9837]=30'd300461633;
array[9838]=30'd432564808;
array[9839]=30'd473528913;
array[9840]=30'd473528913;
array[9841]=30'd488205898;
array[9842]=30'd488205898;
array[9843]=30'd488205898;
array[9844]=30'd473528913;
array[9845]=30'd473528913;
array[9846]=30'd473528913;
array[9847]=30'd458840642;
array[9848]=30'd414803529;
array[9849]=30'd488205898;
array[9850]=30'd488205898;
array[9851]=30'd488205898;
array[9852]=30'd488205898;
array[9853]=30'd488205898;
array[9854]=30'd473528913;
array[9855]=30'd473528913;
array[9856]=30'd458840642;
array[9857]=30'd371776054;
array[9858]=30'd300461633;
array[9859]=30'd453540449;
array[9860]=30'd458840642;
array[9861]=30'd458840642;
array[9862]=30'd315184704;
array[9863]=30'd458840642;
array[9864]=30'd473528913;
array[9865]=30'd352935499;
array[9866]=30'd473528913;
array[9867]=30'd473528913;
array[9868]=30'd473528913;
array[9869]=30'd473528913;
array[9870]=30'd473528913;
array[9871]=30'd458840642;
array[9872]=30'd481853012;
array[9873]=30'd920102487;
array[9874]=30'd920102487;
array[9875]=30'd920102487;
array[9876]=30'd920102487;
array[9877]=30'd920102487;
array[9878]=30'd920102487;
array[9879]=30'd920102487;
array[9880]=30'd920102487;
array[9881]=30'd936883742;
array[9882]=30'd936883742;
array[9883]=30'd875032088;
array[9884]=30'd855119352;
array[9885]=30'd855119352;
array[9886]=30'd855119352;
array[9887]=30'd936883742;
array[9888]=30'd465022394;
array[9889]=30'd478665137;
array[9890]=30'd465022394;
array[9891]=30'd465022394;
array[9892]=30'd465022394;
array[9893]=30'd465022394;
array[9894]=30'd609741283;
array[9895]=30'd915924476;
array[9896]=30'd875032088;
array[9897]=30'd808945195;
array[9898]=30'd756500033;
array[9899]=30'd884420162;
array[9900]=30'd920102487;
array[9901]=30'd920102487;
array[9902]=30'd920102487;
array[9903]=30'd756500033;
array[9904]=30'd860306981;
array[9905]=30'd963075636;
array[9906]=30'd963075636;
array[9907]=30'd963075636;
array[9908]=30'd963075636;
array[9909]=30'd963075636;
array[9910]=30'd963075636;
array[9911]=30'd963075636;
array[9912]=30'd963075636;
array[9913]=30'd963075636;
array[9914]=30'd860306981;
array[9915]=30'd808945195;
array[9916]=30'd920102487;
array[9917]=30'd920102487;
array[9918]=30'd920102487;
array[9919]=30'd920102487;
array[9920]=30'd920102487;
array[9921]=30'd920102487;
array[9922]=30'd920102487;
array[9923]=30'd920102487;
array[9924]=30'd920102487;
array[9925]=30'd920102487;
array[9926]=30'd565736011;
array[9927]=30'd481853012;
array[9928]=30'd473528913;
array[9929]=30'd488205898;
array[9930]=30'd488205898;
array[9931]=30'd488205898;
array[9932]=30'd414803529;
array[9933]=30'd340285012;
array[9934]=30'd381210191;
array[9935]=30'd473528913;
array[9936]=30'd488205898;
array[9937]=30'd488205898;
array[9938]=30'd488205898;
array[9939]=30'd488205898;
array[9940]=30'd488205898;
array[9941]=30'd473528913;
array[9942]=30'd473528913;
array[9943]=30'd414803529;
array[9944]=30'd473528913;
array[9945]=30'd473528913;
array[9946]=30'd488205898;
array[9947]=30'd488205898;
array[9948]=30'd473528913;
array[9949]=30'd488205898;
array[9950]=30'd488205898;
array[9951]=30'd488205898;
array[9952]=30'd473528913;
array[9953]=30'd414803529;
array[9954]=30'd254351946;
array[9955]=30'd458840642;
array[9956]=30'd473528913;
array[9957]=30'd473528913;
array[9958]=30'd458840642;
array[9959]=30'd458840642;
array[9960]=30'd414803529;
array[9961]=30'd414803529;
array[9962]=30'd473528913;
array[9963]=30'd473528913;
array[9964]=30'd473528913;
array[9965]=30'd473528913;
array[9966]=30'd473528913;
array[9967]=30'd473528913;
array[9968]=30'd414803529;
array[9969]=30'd851962439;
array[9970]=30'd920102487;
array[9971]=30'd920102487;
array[9972]=30'd920102487;
array[9973]=30'd920102487;
array[9974]=30'd920102487;
array[9975]=30'd963075636;
array[9976]=30'd915924476;
array[9977]=30'd832058842;
array[9978]=30'd764966339;
array[9979]=30'd778588583;
array[9980]=30'd790145435;
array[9981]=30'd778588583;
array[9982]=30'd764966339;
array[9983]=30'd832058842;
array[9984]=30'd445105582;
array[9985]=30'd489151968;
array[9986]=30'd541577678;
array[9987]=30'd561484289;
array[9988]=30'd650619404;
array[9989]=30'd724009508;
array[9990]=30'd756500033;
array[9991]=30'd808945195;
array[9992]=30'd839339599;
array[9993]=30'd920102487;
array[9994]=30'd920102487;
array[9995]=30'd920102487;
array[9996]=30'd920102487;
array[9997]=30'd920102487;
array[9998]=30'd884420162;
array[9999]=30'd724009508;
array[10000]=30'd778553911;
array[10001]=30'd936883742;
array[10002]=30'd981941808;
array[10003]=30'd963075636;
array[10004]=30'd963075636;
array[10005]=30'd963075636;
array[10006]=30'd963075636;
array[10007]=30'd963075636;
array[10008]=30'd963075636;
array[10009]=30'd860306981;
array[10010]=30'd681011766;
array[10011]=30'd941029952;
array[10012]=30'd920102487;
array[10013]=30'd920102487;
array[10014]=30'd920102487;
array[10015]=30'd920102487;
array[10016]=30'd920102487;
array[10017]=30'd920102487;
array[10018]=30'd920102487;
array[10019]=30'd920102487;
array[10020]=30'd920102487;
array[10021]=30'd650670663;
array[10022]=30'd481853012;
array[10023]=30'd488205898;
array[10024]=30'd488205898;
array[10025]=30'd488205898;
array[10026]=30'd488205898;
array[10027]=30'd458840642;
array[10028]=30'd414803529;
array[10029]=30'd458840642;
array[10030]=30'd352935499;
array[10031]=30'd458840642;
array[10032]=30'd473528913;
array[10033]=30'd473528913;
array[10034]=30'd488205898;
array[10035]=30'd473528913;
array[10036]=30'd473528913;
array[10037]=30'd473528913;
array[10038]=30'd458840642;
array[10039]=30'd414803529;
array[10040]=30'd473528913;
array[10041]=30'd473528913;
array[10042]=30'd488205898;
array[10043]=30'd488205898;
array[10044]=30'd473528913;
array[10045]=30'd488205898;
array[10046]=30'd473528913;
array[10047]=30'd473528913;
array[10048]=30'd458840642;
array[10049]=30'd481853012;
array[10050]=30'd340285012;
array[10051]=30'd481853012;
array[10052]=30'd473528913;
array[10053]=30'd473528913;
array[10054]=30'd473528913;
array[10055]=30'd473528913;
array[10056]=30'd352935499;
array[10057]=30'd473528913;
array[10058]=30'd473528913;
array[10059]=30'd473528913;
array[10060]=30'd473528913;
array[10061]=30'd473528913;
array[10062]=30'd473528913;
array[10063]=30'd473528913;
array[10064]=30'd458840642;
array[10065]=30'd726149706;
array[10066]=30'd920102487;
array[10067]=30'd920102487;
array[10068]=30'd920102487;
array[10069]=30'd920102487;
array[10070]=30'd963075636;
array[10071]=30'd936883742;
array[10072]=30'd785935846;
array[10073]=30'd790145435;
array[10074]=30'd834187654;
array[10075]=30'd854099361;
array[10076]=30'd883468684;
array[10077]=30'd944268729;
array[10078]=30'd854099361;
array[10079]=30'd778588583;
array[10080]=30'd810051001;
array[10081]=30'd896012764;
array[10082]=30'd983039487;
array[10083]=30'd936883742;
array[10084]=30'd936883742;
array[10085]=30'd920102487;
array[10086]=30'd920102487;
array[10087]=30'd920102487;
array[10088]=30'd920102487;
array[10089]=30'd920102487;
array[10090]=30'd920102487;
array[10091]=30'd920102487;
array[10092]=30'd920102487;
array[10093]=30'd884420162;
array[10094]=30'd808945195;
array[10095]=30'd963075636;
array[10096]=30'd936883742;
array[10097]=30'd778553911;
array[10098]=30'd963075636;
array[10099]=30'd963075636;
array[10100]=30'd963075636;
array[10101]=30'd963075636;
array[10102]=30'd963075636;
array[10103]=30'd963075636;
array[10104]=30'd808945195;
array[10105]=30'd793183798;
array[10106]=30'd808945195;
array[10107]=30'd808945195;
array[10108]=30'd963075636;
array[10109]=30'd920102487;
array[10110]=30'd920102487;
array[10111]=30'd920102487;
array[10112]=30'd920102487;
array[10113]=30'd920102487;
array[10114]=30'd920102487;
array[10115]=30'd920102487;
array[10116]=30'd650670663;
array[10117]=30'd481853012;
array[10118]=30'd488205898;
array[10119]=30'd473528913;
array[10120]=30'd473528913;
array[10121]=30'd488205898;
array[10122]=30'd458840642;
array[10123]=30'd414803529;
array[10124]=30'd473528913;
array[10125]=30'd488205898;
array[10126]=30'd473528913;
array[10127]=30'd458840642;
array[10128]=30'd473528913;
array[10129]=30'd488205898;
array[10130]=30'd473528913;
array[10131]=30'd473528913;
array[10132]=30'd473528913;
array[10133]=30'd473528913;
array[10134]=30'd352935499;
array[10135]=30'd458840642;
array[10136]=30'd473528913;
array[10137]=30'd473528913;
array[10138]=30'd473528913;
array[10139]=30'd488205898;
array[10140]=30'd488205898;
array[10141]=30'd473528913;
array[10142]=30'd473528913;
array[10143]=30'd473528913;
array[10144]=30'd543728178;
array[10145]=30'd808945195;
array[10146]=30'd641178184;
array[10147]=30'd650670663;
array[10148]=30'd458840642;
array[10149]=30'd458840642;
array[10150]=30'd473528913;
array[10151]=30'd458840642;
array[10152]=30'd315184704;
array[10153]=30'd458840642;
array[10154]=30'd414803529;
array[10155]=30'd458840642;
array[10156]=30'd473528913;
array[10157]=30'd473528913;
array[10158]=30'd473528913;
array[10159]=30'd473528913;
array[10160]=30'd458840642;
array[10161]=30'd518575683;
array[10162]=30'd920102487;
array[10163]=30'd920102487;
array[10164]=30'd920102487;
array[10165]=30'd963075636;
array[10166]=30'd1002945052;
array[10167]=30'd832058842;
array[10168]=30'd790145435;
array[10169]=30'd914919842;
array[10170]=30'd883468684;
array[10171]=30'd790145435;
array[10172]=30'd854099361;
array[10173]=30'd963129822;
array[10174]=30'd944268729;
array[10175]=30'd778588583;
array[10176]=30'd810051001;
array[10177]=30'd896012764;
array[10178]=30'd963129822;
array[10179]=30'd832058842;
array[10180]=30'd936883742;
array[10181]=30'd920102487;
array[10182]=30'd920102487;
array[10183]=30'd920102487;
array[10184]=30'd920102487;
array[10185]=30'd920102487;
array[10186]=30'd920102487;
array[10187]=30'd920102487;
array[10188]=30'd898096696;
array[10189]=30'd808945195;
array[10190]=30'd1002945052;
array[10191]=30'd1002945052;
array[10192]=30'd936883742;
array[10193]=30'd681011766;
array[10194]=30'd756500033;
array[10195]=30'd860306981;
array[10196]=30'd963075636;
array[10197]=30'd963075636;
array[10198]=30'd884420162;
array[10199]=30'd756500033;
array[10200]=30'd884420162;
array[10201]=30'd963075636;
array[10202]=30'd963075636;
array[10203]=30'd756500033;
array[10204]=30'd884420162;
array[10205]=30'd920102487;
array[10206]=30'd920102487;
array[10207]=30'd920102487;
array[10208]=30'd920102487;
array[10209]=30'd920102487;
array[10210]=30'd920102487;
array[10211]=30'd726149706;
array[10212]=30'd453540449;
array[10213]=30'd488205898;
array[10214]=30'd488205898;
array[10215]=30'd488205898;
array[10216]=30'd473528913;
array[10217]=30'd473528913;
array[10218]=30'd414803529;
array[10219]=30'd473528913;
array[10220]=30'd473528913;
array[10221]=30'd488205898;
array[10222]=30'd488205898;
array[10223]=30'd473528913;
array[10224]=30'd488205898;
array[10225]=30'd488205898;
array[10226]=30'd488205898;
array[10227]=30'd488205898;
array[10228]=30'd352935499;
array[10229]=30'd414803529;
array[10230]=30'd352935499;
array[10231]=30'd473528913;
array[10232]=30'd473528913;
array[10233]=30'd473528913;
array[10234]=30'd473528913;
array[10235]=30'd473528913;
array[10236]=30'd488205898;
array[10237]=30'd488205898;
array[10238]=30'd473528913;
array[10239]=30'd518575683;
array[10240]=30'd851962439;
array[10241]=30'd641178184;
array[10242]=30'd712433198;
array[10243]=30'd641178184;
array[10244]=30'd481853012;
array[10245]=30'd458840642;
array[10246]=30'd458840642;
array[10247]=30'd414803529;
array[10248]=30'd819475993;
array[10249]=30'd898096696;
array[10250]=30'd898096696;
array[10251]=30'd543728178;
array[10252]=30'd458840642;
array[10253]=30'd473528913;
array[10254]=30'd473528913;
array[10255]=30'd473528913;
array[10256]=30'd473528913;
array[10257]=30'd458840642;
array[10258]=30'd726149706;
array[10259]=30'd920102487;
array[10260]=30'd963075636;
array[10261]=30'd963075636;
array[10262]=30'd915924476;
array[10263]=30'd764966339;
array[10264]=30'd854099361;
array[10265]=30'd854099361;
array[10266]=30'd763929993;
array[10267]=30'd763929993;
array[10268]=30'd778588583;
array[10269]=30'd926409165;
array[10270]=30'd979925417;
array[10271]=30'd790145435;
array[10272]=30'd810051001;
array[10273]=30'd926409165;
array[10274]=30'd963129822;
array[10275]=30'd832058842;
array[10276]=30'd915924476;
array[10277]=30'd916923947;
array[10278]=30'd920102487;
array[10279]=30'd920102487;
array[10280]=30'd920102487;
array[10281]=30'd920102487;
array[10282]=30'd920102487;
array[10283]=30'd851962439;
array[10284]=30'd808945195;
array[10285]=30'd1002945052;
array[10286]=30'd1002945052;
array[10287]=30'd963077644;
array[10288]=30'd778553911;
array[10289]=30'd898096696;
array[10290]=30'd920102487;
array[10291]=30'd808945195;
array[10292]=30'd724009508;
array[10293]=30'd556235306;
array[10294]=30'd778553911;
array[10295]=30'd963075636;
array[10296]=30'd963075636;
array[10297]=30'd963075636;
array[10298]=30'd963075636;
array[10299]=30'd941029952;
array[10300]=30'd756500033;
array[10301]=30'd920102487;
array[10302]=30'd920102487;
array[10303]=30'd920102487;
array[10304]=30'd920102487;
array[10305]=30'd920102487;
array[10306]=30'd726149706;
array[10307]=30'd453540449;
array[10308]=30'd518575683;
array[10309]=30'd488205898;
array[10310]=30'd473528913;
array[10311]=30'd488205898;
array[10312]=30'd473528913;
array[10313]=30'd414803529;
array[10314]=30'd458840642;
array[10315]=30'd473528913;
array[10316]=30'd488205898;
array[10317]=30'd488205898;
array[10318]=30'd488205898;
array[10319]=30'd488205898;
array[10320]=30'd488205898;
array[10321]=30'd488205898;
array[10322]=30'd473528913;
array[10323]=30'd473528913;
array[10324]=30'd414803529;
array[10325]=30'd352935499;
array[10326]=30'd458840642;
array[10327]=30'd473528913;
array[10328]=30'd473528913;
array[10329]=30'd473528913;
array[10330]=30'd473528913;
array[10331]=30'd473528913;
array[10332]=30'd488205898;
array[10333]=30'd488205898;
array[10334]=30'd488205898;
array[10335]=30'd518575683;
array[10336]=30'd726149706;
array[10337]=30'd756500033;
array[10338]=30'd793183798;
array[10339]=30'd724009508;
array[10340]=30'd482884128;
array[10341]=30'd494467625;
array[10342]=30'd494467625;
array[10343]=30'd415828509;
array[10344]=30'd808945195;
array[10345]=30'd808945195;
array[10346]=30'd808945195;
array[10347]=30'd586701367;
array[10348]=30'd432564808;
array[10349]=30'd473528913;
array[10350]=30'd473528913;
array[10351]=30'd473528913;
array[10352]=30'd473528913;
array[10353]=30'd473528913;
array[10354]=30'd414803529;
array[10355]=30'd851962439;
array[10356]=30'd963075636;
array[10357]=30'd983039487;
array[10358]=30'd832058842;
array[10359]=30'd790145435;
array[10360]=30'd834187654;
array[10361]=30'd763929993;
array[10362]=30'd790145435;
array[10363]=30'd914919842;
array[10364]=30'd854099361;
array[10365]=30'd914919842;
array[10366]=30'd914919842;
array[10367]=30'd750292390;
array[10368]=30'd852917899;
array[10369]=30'd852917899;
array[10370]=30'd852917899;
array[10371]=30'd852917899;
array[10372]=30'd852917899;
array[10373]=30'd852917899;
array[10374]=30'd852917899;
array[10375]=30'd852917899;
array[10376]=30'd852917899;
array[10377]=30'd852917899;
array[10378]=30'd852917899;
array[10379]=30'd852917899;
array[10380]=30'd852917899;
array[10381]=30'd852917899;
array[10382]=30'd852917899;
array[10383]=30'd852917899;
array[10384]=30'd852917899;
array[10385]=30'd852917899;
array[10386]=30'd852917899;
array[10387]=30'd852917899;
array[10388]=30'd852917899;
array[10389]=30'd852917899;
array[10390]=30'd852917899;
array[10391]=30'd852917899;
array[10392]=30'd852917899;
array[10393]=30'd852917899;
array[10394]=30'd852917899;
array[10395]=30'd873911932;
array[10396]=30'd873911932;
array[10397]=30'd840392271;
array[10398]=30'd910663171;
array[10399]=30'd888658404;
array[10400]=30'd869807552;
array[10401]=30'd832058842;
array[10402]=30'd870795757;
array[10403]=30'd887567935;
array[10404]=30'd852917899;
array[10405]=30'd852917899;
array[10406]=30'd852917899;
array[10407]=30'd852917899;
array[10408]=30'd852917899;
array[10409]=30'd852917899;
array[10410]=30'd852917899;
array[10411]=30'd773214847;
array[10412]=30'd461756049;
array[10413]=30'd461756049;
array[10414]=30'd557159098;
array[10415]=30'd596983478;
array[10416]=30'd596983478;
array[10417]=30'd546644676;
array[10418]=30'd632612564;
array[10419]=30'd632612564;
array[10420]=30'd596983478;
array[10421]=30'd596983478;
array[10422]=30'd632612564;
array[10423]=30'd632612564;
array[10424]=30'd596983478;
array[10425]=30'd653676161;
array[10426]=30'd522581659;
array[10427]=30'd644165300;
array[10428]=30'd650433234;
array[10429]=30'd632612564;
array[10430]=30'd632612564;
array[10431]=30'd650433234;
array[10432]=30'd650433234;
array[10433]=30'd650433234;
array[10434]=30'd632612564;
array[10435]=30'd632612564;
array[10436]=30'd632612564;
array[10437]=30'd596983478;
array[10438]=30'd355833516;
array[10439]=30'd596983478;
array[10440]=30'd644165300;
array[10441]=30'd632612564;
array[10442]=30'd632612564;
array[10443]=30'd632612564;
array[10444]=30'd632612564;
array[10445]=30'd650433234;
array[10446]=30'd644165300;
array[10447]=30'd557159098;
array[10448]=30'd792127082;
array[10449]=30'd792127082;
array[10450]=30'd821480030;
array[10451]=30'd815162003;
array[10452]=30'd815162003;
array[10453]=30'd852917899;
array[10454]=30'd815162003;
array[10455]=30'd852917899;
array[10456]=30'd852917899;
array[10457]=30'd852917899;
array[10458]=30'd852917899;
array[10459]=30'd852917899;
array[10460]=30'd852917899;
array[10461]=30'd852917899;
array[10462]=30'd852917899;
array[10463]=30'd873911932;
array[10464]=30'd852917899;
array[10465]=30'd852917899;
array[10466]=30'd852917899;
array[10467]=30'd852917899;
array[10468]=30'd852917899;
array[10469]=30'd852917899;
array[10470]=30'd852917899;
array[10471]=30'd852917899;
array[10472]=30'd852917899;
array[10473]=30'd852917899;
array[10474]=30'd852917899;
array[10475]=30'd852917899;
array[10476]=30'd852917899;
array[10477]=30'd852917899;
array[10478]=30'd852917899;
array[10479]=30'd852917899;
array[10480]=30'd852917899;
array[10481]=30'd852917899;
array[10482]=30'd852917899;
array[10483]=30'd852917899;
array[10484]=30'd852917899;
array[10485]=30'd852917899;
array[10486]=30'd852917899;
array[10487]=30'd852917899;
array[10488]=30'd852917899;
array[10489]=30'd852917899;
array[10490]=30'd852917899;
array[10491]=30'd852917899;
array[10492]=30'd873911932;
array[10493]=30'd840392271;
array[10494]=30'd916923947;
array[10495]=30'd844591615;
array[10496]=30'd844591615;
array[10497]=30'd862402083;
array[10498]=30'd862402083;
array[10499]=30'd867617357;
array[10500]=30'd852917899;
array[10501]=30'd852917899;
array[10502]=30'd852917899;
array[10503]=30'd852917899;
array[10504]=30'd852917899;
array[10505]=30'd852917899;
array[10506]=30'd852917899;
array[10507]=30'd560346760;
array[10508]=30'd452327079;
array[10509]=30'd609598119;
array[10510]=30'd444947126;
array[10511]=30'd644165300;
array[10512]=30'd515208870;
array[10513]=30'd596983478;
array[10514]=30'd644165300;
array[10515]=30'd644165300;
array[10516]=30'd515208870;
array[10517]=30'd632612564;
array[10518]=30'd650433234;
array[10519]=30'd644165300;
array[10520]=30'd549823127;
array[10521]=30'd821480030;
array[10522]=30'd527847013;
array[10523]=30'd644165300;
array[10524]=30'd632612564;
array[10525]=30'd632612564;
array[10526]=30'd632612564;
array[10527]=30'd650433234;
array[10528]=30'd650433234;
array[10529]=30'd650433234;
array[10530]=30'd632612564;
array[10531]=30'd632612564;
array[10532]=30'd632612564;
array[10533]=30'd644165300;
array[10534]=30'd387282600;
array[10535]=30'd452327079;
array[10536]=30'd644165300;
array[10537]=30'd632612564;
array[10538]=30'd632612564;
array[10539]=30'd632612564;
array[10540]=30'd604303067;
array[10541]=30'd632612564;
array[10542]=30'd632612564;
array[10543]=30'd609598119;
array[10544]=30'd740728401;
array[10545]=30'd887567935;
array[10546]=30'd821480030;
array[10547]=30'd815162003;
array[10548]=30'd815162003;
array[10549]=30'd815162003;
array[10550]=30'd815162003;
array[10551]=30'd852917899;
array[10552]=30'd852917899;
array[10553]=30'd852917899;
array[10554]=30'd852917899;
array[10555]=30'd852917899;
array[10556]=30'd852917899;
array[10557]=30'd873911932;
array[10558]=30'd900139626;
array[10559]=30'd921150041;
array[10560]=30'd852917899;
array[10561]=30'd852917899;
array[10562]=30'd852917899;
array[10563]=30'd852917899;
array[10564]=30'd852917899;
array[10565]=30'd852917899;
array[10566]=30'd852917899;
array[10567]=30'd852917899;
array[10568]=30'd852917899;
array[10569]=30'd852917899;
array[10570]=30'd852917899;
array[10571]=30'd852917899;
array[10572]=30'd852917899;
array[10573]=30'd852917899;
array[10574]=30'd852917899;
array[10575]=30'd852917899;
array[10576]=30'd852917899;
array[10577]=30'd852917899;
array[10578]=30'd852917899;
array[10579]=30'd852917899;
array[10580]=30'd852917899;
array[10581]=30'd852917899;
array[10582]=30'd852917899;
array[10583]=30'd852917899;
array[10584]=30'd852917899;
array[10585]=30'd852917899;
array[10586]=30'd852917899;
array[10587]=30'd852917899;
array[10588]=30'd852917899;
array[10589]=30'd852917899;
array[10590]=30'd867617357;
array[10591]=30'd867617357;
array[10592]=30'd867617357;
array[10593]=30'd867617357;
array[10594]=30'd867617357;
array[10595]=30'd852917899;
array[10596]=30'd852917899;
array[10597]=30'd852917899;
array[10598]=30'd852917899;
array[10599]=30'd852917899;
array[10600]=30'd852917899;
array[10601]=30'd852917899;
array[10602]=30'd773214847;
array[10603]=30'd452327079;
array[10604]=30'd461756049;
array[10605]=30'd609598119;
array[10606]=30'd485848753;
array[10607]=30'd644165300;
array[10608]=30'd485848753;
array[10609]=30'd644165300;
array[10610]=30'd632612564;
array[10611]=30'd644165300;
array[10612]=30'd485848753;
array[10613]=30'd632612564;
array[10614]=30'd650433234;
array[10615]=30'd557159098;
array[10616]=30'd740735615;
array[10617]=30'd804758111;
array[10618]=30'd527847013;
array[10619]=30'd644165300;
array[10620]=30'd632612564;
array[10621]=30'd632612564;
array[10622]=30'd632612564;
array[10623]=30'd650433234;
array[10624]=30'd632612564;
array[10625]=30'd650433234;
array[10626]=30'd632612564;
array[10627]=30'd632612564;
array[10628]=30'd650433234;
array[10629]=30'd632612564;
array[10630]=30'd515208870;
array[10631]=30'd364251806;
array[10632]=30'd644165300;
array[10633]=30'd632612564;
array[10634]=30'd650433234;
array[10635]=30'd632612564;
array[10636]=30'd546644676;
array[10637]=30'd604303067;
array[10638]=30'd632612564;
array[10639]=30'd644165300;
array[10640]=30'd560346760;
array[10641]=30'd821480030;
array[10642]=30'd821480030;
array[10643]=30'd815162003;
array[10644]=30'd815162003;
array[10645]=30'd815162003;
array[10646]=30'd852917899;
array[10647]=30'd852917899;
array[10648]=30'd852917899;
array[10649]=30'd852917899;
array[10650]=30'd852917899;
array[10651]=30'd873911932;
array[10652]=30'd900139626;
array[10653]=30'd959928886;
array[10654]=30'd967280137;
array[10655]=30'd926429685;
array[10656]=30'd852917899;
array[10657]=30'd852917899;
array[10658]=30'd852917899;
array[10659]=30'd852917899;
array[10660]=30'd852917899;
array[10661]=30'd852917899;
array[10662]=30'd852917899;
array[10663]=30'd852917899;
array[10664]=30'd852917899;
array[10665]=30'd852917899;
array[10666]=30'd852917899;
array[10667]=30'd852917899;
array[10668]=30'd852917899;
array[10669]=30'd852917899;
array[10670]=30'd852917899;
array[10671]=30'd852917899;
array[10672]=30'd852917899;
array[10673]=30'd852917899;
array[10674]=30'd852917899;
array[10675]=30'd852917899;
array[10676]=30'd852917899;
array[10677]=30'd852917899;
array[10678]=30'd852917899;
array[10679]=30'd852917899;
array[10680]=30'd852917899;
array[10681]=30'd852917899;
array[10682]=30'd852917899;
array[10683]=30'd852917899;
array[10684]=30'd852917899;
array[10685]=30'd852917899;
array[10686]=30'd852917899;
array[10687]=30'd852917899;
array[10688]=30'd852917899;
array[10689]=30'd852917899;
array[10690]=30'd852917899;
array[10691]=30'd852917899;
array[10692]=30'd852917899;
array[10693]=30'd852917899;
array[10694]=30'd852917899;
array[10695]=30'd852917899;
array[10696]=30'd852917899;
array[10697]=30'd852917899;
array[10698]=30'd653676161;
array[10699]=30'd496374434;
array[10700]=30'd557159098;
array[10701]=30'd557159098;
array[10702]=30'd557159098;
array[10703]=30'd596983478;
array[10704]=30'd515208870;
array[10705]=30'd644165300;
array[10706]=30'd644165300;
array[10707]=30'd485848753;
array[10708]=30'd557159098;
array[10709]=30'd632612564;
array[10710]=30'd644165300;
array[10711]=30'd581297788;
array[10712]=30'd941029952;
array[10713]=30'd840392271;
array[10714]=30'd527847013;
array[10715]=30'd636841618;
array[10716]=30'd546644676;
array[10717]=30'd632612564;
array[10718]=30'd650433234;
array[10719]=30'd604303067;
array[10720]=30'd557159098;
array[10721]=30'd632612564;
array[10722]=30'd632612564;
array[10723]=30'd632612564;
array[10724]=30'd632612564;
array[10725]=30'd632612564;
array[10726]=30'd557159098;
array[10727]=30'd300284569;
array[10728]=30'd609598119;
array[10729]=30'd632612564;
array[10730]=30'd632612564;
array[10731]=30'd632612564;
array[10732]=30'd604303067;
array[10733]=30'd546644676;
array[10734]=30'd632612564;
array[10735]=30'd644165300;
array[10736]=30'd549823127;
array[10737]=30'd740735615;
array[10738]=30'd821480030;
array[10739]=30'd852917899;
array[10740]=30'd852917899;
array[10741]=30'd852917899;
array[10742]=30'd852917899;
array[10743]=30'd852917899;
array[10744]=30'd852917899;
array[10745]=30'd852917899;
array[10746]=30'd852917899;
array[10747]=30'd900139626;
array[10748]=30'd898098744;
array[10749]=30'd910663171;
array[10750]=30'd832058842;
array[10751]=30'd764964292;
array[10752]=30'd852917899;
array[10753]=30'd852917899;
array[10754]=30'd852917899;
array[10755]=30'd852917899;
array[10756]=30'd852917899;
array[10757]=30'd852917899;
array[10758]=30'd852917899;
array[10759]=30'd852917899;
array[10760]=30'd852917899;
array[10761]=30'd852917899;
array[10762]=30'd852917899;
array[10763]=30'd873911932;
array[10764]=30'd873911932;
array[10765]=30'd873911932;
array[10766]=30'd900139626;
array[10767]=30'd867617357;
array[10768]=30'd887567935;
array[10769]=30'd867617357;
array[10770]=30'd867617357;
array[10771]=30'd867617357;
array[10772]=30'd873911932;
array[10773]=30'd900139626;
array[10774]=30'd867617357;
array[10775]=30'd867617357;
array[10776]=30'd852917899;
array[10777]=30'd852917899;
array[10778]=30'd852917899;
array[10779]=30'd852917899;
array[10780]=30'd852917899;
array[10781]=30'd852917899;
array[10782]=30'd852917899;
array[10783]=30'd852917899;
array[10784]=30'd852917899;
array[10785]=30'd852917899;
array[10786]=30'd852917899;
array[10787]=30'd852917899;
array[10788]=30'd852917899;
array[10789]=30'd852917899;
array[10790]=30'd852917899;
array[10791]=30'd852917899;
array[10792]=30'd852917899;
array[10793]=30'd815162003;
array[10794]=30'd496374434;
array[10795]=30'd461756049;
array[10796]=30'd636841618;
array[10797]=30'd515208870;
array[10798]=30'd596983478;
array[10799]=30'd549823127;
array[10800]=30'd557159098;
array[10801]=30'd632612564;
array[10802]=30'd644165300;
array[10803]=30'd496374434;
array[10804]=30'd557159098;
array[10805]=30'd644165300;
array[10806]=30'd609598119;
array[10807]=30'd740728401;
array[10808]=30'd941029952;
array[10809]=30'd867617357;
array[10810]=30'd527847013;
array[10811]=30'd636841618;
array[10812]=30'd444947126;
array[10813]=30'd609598119;
array[10814]=30'd632612564;
array[10815]=30'd644165300;
array[10816]=30'd427157133;
array[10817]=30'd644165300;
array[10818]=30'd650433234;
array[10819]=30'd632612564;
array[10820]=30'd650433234;
array[10821]=30'd596983478;
array[10822]=30'd596983478;
array[10823]=30'd328601227;
array[10824]=30'd522581659;
array[10825]=30'd632612564;
array[10826]=30'd632612564;
array[10827]=30'd632612564;
array[10828]=30'd632612564;
array[10829]=30'd546644676;
array[10830]=30'd644165300;
array[10831]=30'd644165300;
array[10832]=30'd596983478;
array[10833]=30'd710295175;
array[10834]=30'd852917899;
array[10835]=30'd852917899;
array[10836]=30'd852917899;
array[10837]=30'd852917899;
array[10838]=30'd852917899;
array[10839]=30'd852917899;
array[10840]=30'd852917899;
array[10841]=30'd852917899;
array[10842]=30'd852917899;
array[10843]=30'd867617357;
array[10844]=30'd840392271;
array[10845]=30'd778567150;
array[10846]=30'd778567150;
array[10847]=30'd844591615;
array[10848]=30'd852917899;
array[10849]=30'd852917899;
array[10850]=30'd852917899;
array[10851]=30'd852917899;
array[10852]=30'd852917899;
array[10853]=30'd852917899;
array[10854]=30'd852917899;
array[10855]=30'd852917899;
array[10856]=30'd852917899;
array[10857]=30'd852917899;
array[10858]=30'd873911932;
array[10859]=30'd900139626;
array[10860]=30'd921150041;
array[10861]=30'd935829023;
array[10862]=30'd875034136;
array[10863]=30'd855119352;
array[10864]=30'd844591615;
array[10865]=30'd844591615;
array[10866]=30'd844591615;
array[10867]=30'd862402083;
array[10868]=30'd916923947;
array[10869]=30'd959928886;
array[10870]=30'd809995819;
array[10871]=30'd844591615;
array[10872]=30'd867617357;
array[10873]=30'd852917899;
array[10874]=30'd852917899;
array[10875]=30'd852917899;
array[10876]=30'd852917899;
array[10877]=30'd852917899;
array[10878]=30'd852917899;
array[10879]=30'd852917899;
array[10880]=30'd852917899;
array[10881]=30'd852917899;
array[10882]=30'd852917899;
array[10883]=30'd852917899;
array[10884]=30'd852917899;
array[10885]=30'd852917899;
array[10886]=30'd852917899;
array[10887]=30'd852917899;
array[10888]=30'd852917899;
array[10889]=30'd740735615;
array[10890]=30'd496374434;
array[10891]=30'd452327079;
array[10892]=30'd644165300;
array[10893]=30'd444947126;
array[10894]=30'd653646508;
array[10895]=30'd522581659;
array[10896]=30'd596983478;
array[10897]=30'd644165300;
array[10898]=30'd557159098;
array[10899]=30'd604360306;
array[10900]=30'd604360306;
array[10901]=30'd644165300;
array[10902]=30'd549823127;
array[10903]=30'd867617357;
array[10904]=30'd941029952;
array[10905]=30'd887567935;
array[10906]=30'd511088198;
array[10907]=30'd626373227;
array[10908]=30'd626373227;
array[10909]=30'd581297788;
array[10910]=30'd644165300;
array[10911]=30'd644165300;
array[10912]=30'd496374434;
array[10913]=30'd549823127;
array[10914]=30'd644165300;
array[10915]=30'd632612564;
array[10916]=30'd632612564;
array[10917]=30'd485848753;
array[10918]=30'd596983478;
array[10919]=30'd328601227;
array[10920]=30'd427157133;
array[10921]=30'd644165300;
array[10922]=30'd632612564;
array[10923]=30'd650433234;
array[10924]=30'd632612564;
array[10925]=30'd596983478;
array[10926]=30'd546644676;
array[10927]=30'd644165300;
array[10928]=30'd644165300;
array[10929]=30'd609598119;
array[10930]=30'd852917899;
array[10931]=30'd852917899;
array[10932]=30'd815162003;
array[10933]=30'd852917899;
array[10934]=30'd852917899;
array[10935]=30'd852917899;
array[10936]=30'd852917899;
array[10937]=30'd852917899;
array[10938]=30'd852917899;
array[10939]=30'd852917899;
array[10940]=30'd873911932;
array[10941]=30'd840392271;
array[10942]=30'd840392271;
array[10943]=30'd887567935;
array[10944]=30'd852917899;
array[10945]=30'd852917899;
array[10946]=30'd852917899;
array[10947]=30'd852917899;
array[10948]=30'd852917899;
array[10949]=30'd852917899;
array[10950]=30'd852917899;
array[10951]=30'd852917899;
array[10952]=30'd852917899;
array[10953]=30'd873911932;
array[10954]=30'd900139626;
array[10955]=30'd959928886;
array[10956]=30'd950544914;
array[10957]=30'd832058842;
array[10958]=30'd782796193;
array[10959]=30'd782796193;
array[10960]=30'd768126344;
array[10961]=30'd782796193;
array[10962]=30'd764964292;
array[10963]=30'd752351692;
array[10964]=30'd844591615;
array[10965]=30'd967280137;
array[10966]=30'd832058842;
array[10967]=30'd778567150;
array[10968]=30'd862402083;
array[10969]=30'd867617357;
array[10970]=30'd852917899;
array[10971]=30'd852917899;
array[10972]=30'd852917899;
array[10973]=30'd852917899;
array[10974]=30'd852917899;
array[10975]=30'd852917899;
array[10976]=30'd852917899;
array[10977]=30'd852917899;
array[10978]=30'd852917899;
array[10979]=30'd852917899;
array[10980]=30'd852917899;
array[10981]=30'd852917899;
array[10982]=30'd852917899;
array[10983]=30'd852917899;
array[10984]=30'd852917899;
array[10985]=30'd625391195;
array[10986]=30'd560346760;
array[10987]=30'd522581659;
array[10988]=30'd644165300;
array[10989]=30'd444947126;
array[10990]=30'd644165300;
array[10991]=30'd427157133;
array[10992]=30'd644165300;
array[10993]=30'd644165300;
array[10994]=30'd522581659;
array[10995]=30'd740728401;
array[10996]=30'd604360306;
array[10997]=30'd644165300;
array[10998]=30'd653676161;
array[10999]=30'd941029952;
array[11000]=30'd941029952;
array[11001]=30'd941029952;
array[11002]=30'd553016910;
array[11003]=30'd604360306;
array[11004]=30'd757545539;
array[11005]=30'd527847013;
array[11006]=30'd636841618;
array[11007]=30'd644165300;
array[11008]=30'd626373227;
array[11009]=30'd593947240;
array[11010]=30'd636841618;
array[11011]=30'd644165300;
array[11012]=30'd604303067;
array[11013]=30'd444947126;
array[11014]=30'd557159098;
array[11015]=30'd364251806;
array[11016]=30'd404111966;
array[11017]=30'd636841618;
array[11018]=30'd632612564;
array[11019]=30'd632612564;
array[11020]=30'd632612564;
array[11021]=30'd604303067;
array[11022]=30'd515208870;
array[11023]=30'd632612564;
array[11024]=30'd644165300;
array[11025]=30'd549823127;
array[11026]=30'd852917899;
array[11027]=30'd852917899;
array[11028]=30'd852917899;
array[11029]=30'd852917899;
array[11030]=30'd852917899;
array[11031]=30'd852917899;
array[11032]=30'd852917899;
array[11033]=30'd852917899;
array[11034]=30'd852917899;
array[11035]=30'd852917899;
array[11036]=30'd852917899;
array[11037]=30'd852917899;
array[11038]=30'd852917899;
array[11039]=30'd921150041;
array[11040]=30'd852917899;
array[11041]=30'd852917899;
array[11042]=30'd852917899;
array[11043]=30'd852917899;
array[11044]=30'd852917899;
array[11045]=30'd852917899;
array[11046]=30'd852917899;
array[11047]=30'd873911932;
array[11048]=30'd873911932;
array[11049]=30'd873911932;
array[11050]=30'd941029952;
array[11051]=30'd950544914;
array[11052]=30'd832058842;
array[11053]=30'd782796193;
array[11054]=30'd885566856;
array[11055]=30'd885566856;
array[11056]=30'd782796193;
array[11057]=30'd906527146;
array[11058]=30'd945318330;
array[11059]=30'd764964292;
array[11060]=30'd820487650;
array[11061]=30'd910663171;
array[11062]=30'd967280137;
array[11063]=30'd794289609;
array[11064]=30'd820487650;
array[11065]=30'd867617357;
array[11066]=30'd852917899;
array[11067]=30'd852917899;
array[11068]=30'd852917899;
array[11069]=30'd852917899;
array[11070]=30'd852917899;
array[11071]=30'd852917899;
array[11072]=30'd852917899;
array[11073]=30'd852917899;
array[11074]=30'd852917899;
array[11075]=30'd852917899;
array[11076]=30'd852917899;
array[11077]=30'd852917899;
array[11078]=30'd852917899;
array[11079]=30'd852917899;
array[11080]=30'd867617357;
array[11081]=30'd527847013;
array[11082]=30'd560346760;
array[11083]=30'd549823127;
array[11084]=30'd644165300;
array[11085]=30'd452327079;
array[11086]=30'd596983478;
array[11087]=30'd364251806;
array[11088]=30'd636841618;
array[11089]=30'd609598119;
array[11090]=30'd593947240;
array[11091]=30'd794232376;
array[11092]=30'd581297788;
array[11093]=30'd609598119;
array[11094]=30'd757545539;
array[11095]=30'd959928886;
array[11096]=30'd941029952;
array[11097]=30'd941029952;
array[11098]=30'd666281541;
array[11099]=30'd593947240;
array[11100]=30'd821480030;
array[11101]=30'd757545539;
array[11102]=30'd581297788;
array[11103]=30'd644165300;
array[11104]=30'd571937394;
array[11105]=30'd794232376;
array[11106]=30'd581297788;
array[11107]=30'd644165300;
array[11108]=30'd644165300;
array[11109]=30'd515208870;
array[11110]=30'd496374434;
array[11111]=30'd427157133;
array[11112]=30'd351684214;
array[11113]=30'd636841618;
array[11114]=30'd632612564;
array[11115]=30'd632612564;
array[11116]=30'd632612564;
array[11117]=30'd604303067;
array[11118]=30'd515208870;
array[11119]=30'd632612564;
array[11120]=30'd632612564;
array[11121]=30'd549823127;
array[11122]=30'd815162003;
array[11123]=30'd852917899;
array[11124]=30'd852917899;
array[11125]=30'd815162003;
array[11126]=30'd852917899;
array[11127]=30'd852917899;
array[11128]=30'd852917899;
array[11129]=30'd852917899;
array[11130]=30'd852917899;
array[11131]=30'd852917899;
array[11132]=30'd852917899;
array[11133]=30'd852917899;
array[11134]=30'd852917899;
array[11135]=30'd887567935;
array[11136]=30'd852917899;
array[11137]=30'd852917899;
array[11138]=30'd852917899;
array[11139]=30'd852917899;
array[11140]=30'd852917899;
array[11141]=30'd852917899;
array[11142]=30'd852917899;
array[11143]=30'd873911932;
array[11144]=30'd873911932;
array[11145]=30'd921150041;
array[11146]=30'd950544914;
array[11147]=30'd832058842;
array[11148]=30'd782796193;
array[11149]=30'd885566856;
array[11150]=30'd833137031;
array[11151]=30'd768126344;
array[11152]=30'd782796193;
array[11153]=30'd869807552;
array[11154]=30'd1000883648;
array[11155]=30'd764964292;
array[11156]=30'd820487650;
array[11157]=30'd890710541;
array[11158]=30'd1004004888;
array[11159]=30'd832058842;
array[11160]=30'd794289609;
array[11161]=30'd862402083;
array[11162]=30'd873911932;
array[11163]=30'd852917899;
array[11164]=30'd852917899;
array[11165]=30'd852917899;
array[11166]=30'd852917899;
array[11167]=30'd852917899;
array[11168]=30'd852917899;
array[11169]=30'd852917899;
array[11170]=30'd852917899;
array[11171]=30'd852917899;
array[11172]=30'd852917899;
array[11173]=30'd852917899;
array[11174]=30'd852917899;
array[11175]=30'd852917899;
array[11176]=30'd821480030;
array[11177]=30'd503733877;
array[11178]=30'd549823127;
array[11179]=30'd549823127;
array[11180]=30'd609598119;
array[11181]=30'd364251806;
array[11182]=30'd549823127;
array[11183]=30'd433483392;
array[11184]=30'd636841618;
array[11185]=30'd609598119;
array[11186]=30'd709314133;
array[11187]=30'd794232376;
array[11188]=30'd527847013;
array[11189]=30'd581297788;
array[11190]=30'd821480030;
array[11191]=30'd959928886;
array[11192]=30'd959928886;
array[11193]=30'd941029952;
array[11194]=30'd794232376;
array[11195]=30'd511088198;
array[11196]=30'd794232376;
array[11197]=30'd916923947;
array[11198]=30'd527847013;
array[11199]=30'd636841618;
array[11200]=30'd503733877;
array[11201]=30'd887567935;
array[11202]=30'd527847013;
array[11203]=30'd636841618;
array[11204]=30'd644165300;
array[11205]=30'd581297788;
array[11206]=30'd503733877;
array[11207]=30'd593947240;
array[11208]=30'd482780758;
array[11209]=30'd636841618;
array[11210]=30'd632612564;
array[11211]=30'd632612564;
array[11212]=30'd632612564;
array[11213]=30'd604303067;
array[11214]=30'd546644676;
array[11215]=30'd644165300;
array[11216]=30'd632612564;
array[11217]=30'd557159098;
array[11218]=30'd815162003;
array[11219]=30'd852917899;
array[11220]=30'd852917899;
array[11221]=30'd815162003;
array[11222]=30'd852917899;
array[11223]=30'd852917899;
array[11224]=30'd852917899;
array[11225]=30'd852917899;
array[11226]=30'd852917899;
array[11227]=30'd852917899;
array[11228]=30'd852917899;
array[11229]=30'd852917899;
array[11230]=30'd852917899;
array[11231]=30'd867617357;
array[11232]=30'd852917899;
array[11233]=30'd852917899;
array[11234]=30'd852917899;
array[11235]=30'd852917899;
array[11236]=30'd852917899;
array[11237]=30'd852917899;
array[11238]=30'd873911932;
array[11239]=30'd873911932;
array[11240]=30'd900139626;
array[11241]=30'd959928886;
array[11242]=30'd888658404;
array[11243]=30'd782796193;
array[11244]=30'd833137031;
array[11245]=30'd768126344;
array[11246]=30'd768126344;
array[11247]=30'd849905057;
array[11248]=30'd811098555;
array[11249]=30'd869807552;
array[11250]=30'd979923369;
array[11251]=30'd764964292;
array[11252]=30'd820487650;
array[11253]=30'd935829023;
array[11254]=30'd1004004888;
array[11255]=30'd832058842;
array[11256]=30'd794289609;
array[11257]=30'd862402083;
array[11258]=30'd867617357;
array[11259]=30'd852917899;
array[11260]=30'd852917899;
array[11261]=30'd852917899;
array[11262]=30'd852917899;
array[11263]=30'd852917899;
array[11264]=30'd852917899;
array[11265]=30'd852917899;
array[11266]=30'd852917899;
array[11267]=30'd852917899;
array[11268]=30'd852917899;
array[11269]=30'd852917899;
array[11270]=30'd852917899;
array[11271]=30'd852917899;
array[11272]=30'd773214847;
array[11273]=30'd560346760;
array[11274]=30'd557159098;
array[11275]=30'd549823127;
array[11276]=30'd609598119;
array[11277]=30'd328601227;
array[11278]=30'd503733877;
array[11279]=30'd666281541;
array[11280]=30'd581297788;
array[11281]=30'd527847013;
array[11282]=30'd666281541;
array[11283]=30'd794232376;
array[11284]=30'd511088198;
array[11285]=30'd503733877;
array[11286]=30'd794232376;
array[11287]=30'd959928886;
array[11288]=30'd959928886;
array[11289]=30'd959928886;
array[11290]=30'd916923947;
array[11291]=30'd482780758;
array[11292]=30'd642228804;
array[11293]=30'd679964212;
array[11294]=30'd713478705;
array[11295]=30'd560346760;
array[11296]=30'd503733877;
array[11297]=30'd666281541;
array[11298]=30'd625391195;
array[11299]=30'd581297788;
array[11300]=30'd636841618;
array[11301]=30'd593947240;
array[11302]=30'd593947240;
array[11303]=30'd595020337;
array[11304]=30'd666281541;
array[11305]=30'd626373227;
array[11306]=30'd644165300;
array[11307]=30'd596983478;
array[11308]=30'd604303067;
array[11309]=30'd604303067;
array[11310]=30'd546644676;
array[11311]=30'd596983478;
array[11312]=30'd632612564;
array[11313]=30'd557159098;
array[11314]=30'd773214847;
array[11315]=30'd852917899;
array[11316]=30'd852917899;
array[11317]=30'd852917899;
array[11318]=30'd852917899;
array[11319]=30'd852917899;
array[11320]=30'd852917899;
array[11321]=30'd852917899;
array[11322]=30'd852917899;
array[11323]=30'd852917899;
array[11324]=30'd852917899;
array[11325]=30'd852917899;
array[11326]=30'd852917899;
array[11327]=30'd852917899;
array[11328]=30'd852917899;
array[11329]=30'd852917899;
array[11330]=30'd852917899;
array[11331]=30'd852917899;
array[11332]=30'd852917899;
array[11333]=30'd852917899;
array[11334]=30'd873911932;
array[11335]=30'd873911932;
array[11336]=30'd900139626;
array[11337]=30'd959928886;
array[11338]=30'd832058842;
array[11339]=30'd811098555;
array[11340]=30'd849905057;
array[11341]=30'd750292390;
array[11342]=30'd849905057;
array[11343]=30'd945318330;
array[11344]=30'd906527146;
array[11345]=30'd906527146;
array[11346]=30'd869807552;
array[11347]=30'd764964292;
array[11348]=30'd870795757;
array[11349]=30'd987238908;
array[11350]=30'd926429685;
array[11351]=30'd764964292;
array[11352]=30'd820487650;
array[11353]=30'd867617357;
array[11354]=30'd852917899;
array[11355]=30'd852917899;
array[11356]=30'd852917899;
array[11357]=30'd852917899;
array[11358]=30'd852917899;
array[11359]=30'd852917899;
array[11360]=30'd852917899;
array[11361]=30'd852917899;
array[11362]=30'd852917899;
array[11363]=30'd852917899;
array[11364]=30'd852917899;
array[11365]=30'd852917899;
array[11366]=30'd852917899;
array[11367]=30'd852917899;
array[11368]=30'd710295175;
array[11369]=30'd604360306;
array[11370]=30'd609598119;
array[11371]=30'd496374434;
array[11372]=30'd557159098;
array[11373]=30'd503733877;
array[11374]=30'd482780758;
array[11375]=30'd794232376;
array[11376]=30'd482780758;
array[11377]=30'd553016910;
array[11378]=30'd941029952;
array[11379]=30'd959928886;
array[11380]=30'd713478705;
array[11381]=30'd511088198;
array[11382]=30'd941029952;
array[11383]=30'd959928886;
array[11384]=30'd959928886;
array[11385]=30'd959928886;
array[11386]=30'd959928886;
array[11387]=30'd757545539;
array[11388]=30'd679964212;
array[11389]=30'd959928886;
array[11390]=30'd941029952;
array[11391]=30'd666281541;
array[11392]=30'd553016910;
array[11393]=30'd916923947;
array[11394]=30'd862402083;
array[11395]=30'd527847013;
array[11396]=30'd626373227;
array[11397]=30'd679964212;
array[11398]=30'd666281541;
array[11399]=30'd679964212;
array[11400]=30'd757545539;
array[11401]=30'd581297788;
array[11402]=30'd644165300;
array[11403]=30'd596983478;
array[11404]=30'd604303067;
array[11405]=30'd604303067;
array[11406]=30'd596983478;
array[11407]=30'd546644676;
array[11408]=30'd632612564;
array[11409]=30'd596983478;
array[11410]=30'd710295175;
array[11411]=30'd852917899;
array[11412]=30'd852917899;
array[11413]=30'd852917899;
array[11414]=30'd852917899;
array[11415]=30'd852917899;
array[11416]=30'd852917899;
array[11417]=30'd852917899;
array[11418]=30'd852917899;
array[11419]=30'd852917899;
array[11420]=30'd852917899;
array[11421]=30'd852917899;
array[11422]=30'd852917899;
array[11423]=30'd852917899;
array[11424]=30'd852917899;
array[11425]=30'd852917899;
array[11426]=30'd852917899;
array[11427]=30'd852917899;
array[11428]=30'd852917899;
array[11429]=30'd852917899;
array[11430]=30'd873911932;
array[11431]=30'd873911932;
array[11432]=30'd900139626;
array[11433]=30'd959928886;
array[11434]=30'd832058842;
array[11435]=30'd811098555;
array[11436]=30'd906527146;
array[11437]=30'd782796193;
array[11438]=30'd849905057;
array[11439]=30'd945318330;
array[11440]=30'd869807552;
array[11441]=30'd764964292;
array[11442]=30'd764964292;
array[11443]=30'd832058842;
array[11444]=30'd967280137;
array[11445]=30'd987238908;
array[11446]=30'd832058842;
array[11447]=30'd794289609;
array[11448]=30'd844591615;
array[11449]=30'd867617357;
array[11450]=30'd873911932;
array[11451]=30'd852917899;
array[11452]=30'd852917899;
array[11453]=30'd852917899;
array[11454]=30'd852917899;
array[11455]=30'd852917899;
array[11456]=30'd852917899;
array[11457]=30'd852917899;
array[11458]=30'd852917899;
array[11459]=30'd852917899;
array[11460]=30'd852917899;
array[11461]=30'd852917899;
array[11462]=30'd852917899;
array[11463]=30'd873911932;
array[11464]=30'd625391195;
array[11465]=30'd636841618;
array[11466]=30'd644165300;
array[11467]=30'd444947126;
array[11468]=30'd549823127;
array[11469]=30'd709314133;
array[11470]=30'd417793613;
array[11471]=30'd713478705;
array[11472]=30'd583423551;
array[11473]=30'd553016910;
array[11474]=30'd959928886;
array[11475]=30'd959928886;
array[11476]=30'd887567935;
array[11477]=30'd573005379;
array[11478]=30'd959928886;
array[11479]=30'd959928886;
array[11480]=30'd959928886;
array[11481]=30'd959928886;
array[11482]=30'd959928886;
array[11483]=30'd941029952;
array[11484]=30'd794232376;
array[11485]=30'd985089582;
array[11486]=30'd959928886;
array[11487]=30'd887567935;
array[11488]=30'd528975414;
array[11489]=30'd916923947;
array[11490]=30'd959928886;
array[11491]=30'd713478705;
array[11492]=30'd482780758;
array[11493]=30'd757545539;
array[11494]=30'd721911330;
array[11495]=30'd757545539;
array[11496]=30'd757545539;
array[11497]=30'd482780758;
array[11498]=30'd636841618;
array[11499]=30'd557159098;
array[11500]=30'd596983478;
array[11501]=30'd632612564;
array[11502]=30'd596983478;
array[11503]=30'd546644676;
array[11504]=30'd632612564;
array[11505]=30'd596983478;
array[11506]=30'd710295175;
array[11507]=30'd852917899;
array[11508]=30'd852917899;
array[11509]=30'd852917899;
array[11510]=30'd852917899;
array[11511]=30'd852917899;
array[11512]=30'd852917899;
array[11513]=30'd852917899;
array[11514]=30'd852917899;
array[11515]=30'd852917899;
array[11516]=30'd852917899;
array[11517]=30'd852917899;
array[11518]=30'd852917899;
array[11519]=30'd852917899;
array[11520]=30'd852917899;
array[11521]=30'd852917899;
array[11522]=30'd852917899;
array[11523]=30'd852917899;
array[11524]=30'd852917899;
array[11525]=30'd873911932;
array[11526]=30'd873911932;
array[11527]=30'd873911932;
array[11528]=30'd900139626;
array[11529]=30'd959928886;
array[11530]=30'd855119352;
array[11531]=30'd764964292;
array[11532]=30'd904416730;
array[11533]=30'd849905057;
array[11534]=30'd764964292;
array[11535]=30'd750292390;
array[11536]=30'd764964292;
array[11537]=30'd794289609;
array[11538]=30'd855119352;
array[11539]=30'd910663171;
array[11540]=30'd1004004888;
array[11541]=30'd888658404;
array[11542]=30'd752351692;
array[11543]=30'd844591615;
array[11544]=30'd862402083;
array[11545]=30'd873911932;
array[11546]=30'd873911932;
array[11547]=30'd852917899;
array[11548]=30'd852917899;
array[11549]=30'd852917899;
array[11550]=30'd852917899;
array[11551]=30'd852917899;
array[11552]=30'd852917899;
array[11553]=30'd852917899;
array[11554]=30'd852917899;
array[11555]=30'd852917899;
array[11556]=30'd852917899;
array[11557]=30'd852917899;
array[11558]=30'd852917899;
array[11559]=30'd852917899;
array[11560]=30'd593947240;
array[11561]=30'd636841618;
array[11562]=30'd644165300;
array[11563]=30'd515208870;
array[11564]=30'd522581659;
array[11565]=30'd757545539;
array[11566]=30'd472349226;
array[11567]=30'd941029952;
array[11568]=30'd862402083;
array[11569]=30'd573005379;
array[11570]=30'd959928886;
array[11571]=30'd959928886;
array[11572]=30'd959928886;
array[11573]=30'd916923947;
array[11574]=30'd959928886;
array[11575]=30'd959928886;
array[11576]=30'd959928886;
array[11577]=30'd959928886;
array[11578]=30'd959928886;
array[11579]=30'd959928886;
array[11580]=30'd959928886;
array[11581]=30'd959928886;
array[11582]=30'd959928886;
array[11583]=30'd959928886;
array[11584]=30'd887567935;
array[11585]=30'd941029952;
array[11586]=30'd959928886;
array[11587]=30'd887567935;
array[11588]=30'd511088198;
array[11589]=30'd862402083;
array[11590]=30'd595020337;
array[11591]=30'd809995819;
array[11592]=30'd419882502;
array[11593]=30'd472349226;
array[11594]=30'd453416554;
array[11595]=30'd522581659;
array[11596]=30'd596983478;
array[11597]=30'd632612564;
array[11598]=30'd644165300;
array[11599]=30'd546644676;
array[11600]=30'd650433234;
array[11601]=30'd596983478;
array[11602]=30'd740735615;
array[11603]=30'd852917899;
array[11604]=30'd852917899;
array[11605]=30'd852917899;
array[11606]=30'd852917899;
array[11607]=30'd852917899;
array[11608]=30'd852917899;
array[11609]=30'd852917899;
array[11610]=30'd852917899;
array[11611]=30'd852917899;
array[11612]=30'd852917899;
array[11613]=30'd852917899;
array[11614]=30'd852917899;
array[11615]=30'd852917899;
array[11616]=30'd852917899;
array[11617]=30'd852917899;
array[11618]=30'd852917899;
array[11619]=30'd852917899;
array[11620]=30'd873911932;
array[11621]=30'd873911932;
array[11622]=30'd873911932;
array[11623]=30'd873911932;
array[11624]=30'd873911932;
array[11625]=30'd898098744;
array[11626]=30'd926429685;
array[11627]=30'd764964292;
array[11628]=30'd811098555;
array[11629]=30'd888658404;
array[11630]=30'd778567150;
array[11631]=30'd794289609;
array[11632]=30'd820487650;
array[11633]=30'd855119352;
array[11634]=30'd898098744;
array[11635]=30'd1004004888;
array[11636]=30'd926429685;
array[11637]=30'd794289609;
array[11638]=30'd820487650;
array[11639]=30'd862402083;
array[11640]=30'd867617357;
array[11641]=30'd852917899;
array[11642]=30'd852917899;
array[11643]=30'd852917899;
array[11644]=30'd852917899;
array[11645]=30'd852917899;
array[11646]=30'd852917899;
array[11647]=30'd852917899;
array[11648]=30'd852917899;
array[11649]=30'd852917899;
array[11650]=30'd852917899;
array[11651]=30'd852917899;
array[11652]=30'd852917899;
array[11653]=30'd852917899;
array[11654]=30'd852917899;
array[11655]=30'd852917899;
array[11656]=30'd571937394;
array[11657]=30'd636841618;
array[11658]=30'd644165300;
array[11659]=30'd596983478;
array[11660]=30'd397801110;
array[11661]=30'd757545539;
array[11662]=30'd862402083;
array[11663]=30'd959928886;
array[11664]=30'd959928886;
array[11665]=30'd887567935;
array[11666]=30'd959928886;
array[11667]=30'd959928886;
array[11668]=30'd959928886;
array[11669]=30'd959928886;
array[11670]=30'd959928886;
array[11671]=30'd959928886;
array[11672]=30'd959928886;
array[11673]=30'd959928886;
array[11674]=30'd959928886;
array[11675]=30'd959928886;
array[11676]=30'd959928886;
array[11677]=30'd959928886;
array[11678]=30'd959928886;
array[11679]=30'd959928886;
array[11680]=30'd959928886;
array[11681]=30'd959928886;
array[11682]=30'd959928886;
array[11683]=30'd959928886;
array[11684]=30'd916923947;
array[11685]=30'd959928886;
array[11686]=30'd862402083;
array[11687]=30'd809995819;
array[11688]=30'd651672075;
array[11689]=30'd820487650;
array[11690]=30'd455516734;
array[11691]=30'd486913656;
array[11692]=30'd596983478;
array[11693]=30'd632612564;
array[11694]=30'd632612564;
array[11695]=30'd546644676;
array[11696]=30'd632612564;
array[11697]=30'd557159098;
array[11698]=30'd773214847;
array[11699]=30'd852917899;
array[11700]=30'd852917899;
array[11701]=30'd852917899;
array[11702]=30'd852917899;
array[11703]=30'd852917899;
array[11704]=30'd852917899;
array[11705]=30'd852917899;
array[11706]=30'd852917899;
array[11707]=30'd852917899;
array[11708]=30'd852917899;
array[11709]=30'd852917899;
array[11710]=30'd852917899;
array[11711]=30'd852917899;
array[11712]=30'd852917899;
array[11713]=30'd852917899;
array[11714]=30'd852917899;
array[11715]=30'd852917899;
array[11716]=30'd852917899;
array[11717]=30'd873911932;
array[11718]=30'd873911932;
array[11719]=30'd873911932;
array[11720]=30'd873911932;
array[11721]=30'd900139626;
array[11722]=30'd935829023;
array[11723]=30'd832058842;
array[11724]=30'd764964292;
array[11725]=30'd832058842;
array[11726]=30'd910663171;
array[11727]=30'd910663171;
array[11728]=30'd910663171;
array[11729]=30'd935829023;
array[11730]=30'd926429685;
array[11731]=30'd855119352;
array[11732]=30'd764964292;
array[11733]=30'd794289609;
array[11734]=30'd862402083;
array[11735]=30'd867617357;
array[11736]=30'd852917899;
array[11737]=30'd852917899;
array[11738]=30'd873911932;
array[11739]=30'd873911932;
array[11740]=30'd852917899;
array[11741]=30'd852917899;
array[11742]=30'd852917899;
array[11743]=30'd852917899;
array[11744]=30'd852917899;
array[11745]=30'd852917899;
array[11746]=30'd852917899;
array[11747]=30'd852917899;
array[11748]=30'd852917899;
array[11749]=30'd852917899;
array[11750]=30'd873911932;
array[11751]=30'd852917899;
array[11752]=30'd560346760;
array[11753]=30'd636841618;
array[11754]=30'd644165300;
array[11755]=30'd596983478;
array[11756]=30'd560346760;
array[11757]=30'd757545539;
array[11758]=30'd959928886;
array[11759]=30'd959928886;
array[11760]=30'd959928886;
array[11761]=30'd959928886;
array[11762]=30'd887567935;
array[11763]=30'd862402083;
array[11764]=30'd887567935;
array[11765]=30'd959928886;
array[11766]=30'd959928886;
array[11767]=30'd959928886;
array[11768]=30'd959928886;
array[11769]=30'd959928886;
array[11770]=30'd959928886;
array[11771]=30'd959928886;
array[11772]=30'd959928886;
array[11773]=30'd959928886;
array[11774]=30'd959928886;
array[11775]=30'd959928886;
array[11776]=30'd959928886;
array[11777]=30'd959928886;
array[11778]=30'd959928886;
array[11779]=30'd959928886;
array[11780]=30'd959928886;
array[11781]=30'd959928886;
array[11782]=30'd959928886;
array[11783]=30'd875034136;
array[11784]=30'd651672075;
array[11785]=30'd778567150;
array[11786]=30'd511088198;
array[11787]=30'd486913656;
array[11788]=30'd609598119;
array[11789]=30'd632612564;
array[11790]=30'd604303067;
array[11791]=30'd546644676;
array[11792]=30'd632612564;
array[11793]=30'd557159098;
array[11794]=30'd815162003;
array[11795]=30'd852917899;
array[11796]=30'd852917899;
array[11797]=30'd852917899;
array[11798]=30'd852917899;
array[11799]=30'd852917899;
array[11800]=30'd852917899;
array[11801]=30'd852917899;
array[11802]=30'd852917899;
array[11803]=30'd852917899;
array[11804]=30'd852917899;
array[11805]=30'd852917899;
array[11806]=30'd852917899;
array[11807]=30'd852917899;
array[11808]=30'd852917899;
array[11809]=30'd852917899;
array[11810]=30'd852917899;
array[11811]=30'd873911932;
array[11812]=30'd873911932;
array[11813]=30'd873911932;
array[11814]=30'd873911932;
array[11815]=30'd873911932;
array[11816]=30'd873911932;
array[11817]=30'd873911932;
array[11818]=30'd898098744;
array[11819]=30'd898098744;
array[11820]=30'd785935846;
array[11821]=30'd764964292;
array[11822]=30'd832058842;
array[11823]=30'd832058842;
array[11824]=30'd832058842;
array[11825]=30'd811098555;
array[11826]=30'd764964292;
array[11827]=30'd794289609;
array[11828]=30'd820487650;
array[11829]=30'd844591615;
array[11830]=30'd867617357;
array[11831]=30'd873911932;
array[11832]=30'd852917899;
array[11833]=30'd852917899;
array[11834]=30'd852917899;
array[11835]=30'd873911932;
array[11836]=30'd852917899;
array[11837]=30'd852917899;
array[11838]=30'd852917899;
array[11839]=30'd852917899;
array[11840]=30'd852917899;
array[11841]=30'd852917899;
array[11842]=30'd873911932;
array[11843]=30'd873911932;
array[11844]=30'd852917899;
array[11845]=30'd852917899;
array[11846]=30'd852917899;
array[11847]=30'd852917899;
array[11848]=30'd581297788;
array[11849]=30'd636841618;
array[11850]=30'd644165300;
array[11851]=30'd515208870;
array[11852]=30'd609598119;
array[11853]=30'd757545539;
array[11854]=30'd959928886;
array[11855]=30'd959928886;
array[11856]=30'd862402083;
array[11857]=30'd721911330;
array[11858]=30'd757545539;
array[11859]=30'd862402083;
array[11860]=30'd809995819;
array[11861]=30'd809995819;
array[11862]=30'd959928886;
array[11863]=30'd959928886;
array[11864]=30'd959928886;
array[11865]=30'd959928886;
array[11866]=30'd959928886;
array[11867]=30'd959928886;
array[11868]=30'd959928886;
array[11869]=30'd916923947;
array[11870]=30'd809995819;
array[11871]=30'd721911330;
array[11872]=30'd721911330;
array[11873]=30'd757545539;
array[11874]=30'd916923947;
array[11875]=30'd959928886;
array[11876]=30'd959928886;
array[11877]=30'd959928886;
array[11878]=30'd959928886;
array[11879]=30'd862402083;
array[11880]=30'd501707283;
array[11881]=30'd472349226;
array[11882]=30'd553016910;
array[11883]=30'd486913656;
array[11884]=30'd644165300;
array[11885]=30'd632612564;
array[11886]=30'd644165300;
array[11887]=30'd557159098;
array[11888]=30'd632612564;
array[11889]=30'd549823127;
array[11890]=30'd815162003;
array[11891]=30'd852917899;
array[11892]=30'd852917899;
array[11893]=30'd852917899;
array[11894]=30'd852917899;
array[11895]=30'd852917899;
array[11896]=30'd852917899;
array[11897]=30'd852917899;
array[11898]=30'd852917899;
array[11899]=30'd852917899;
array[11900]=30'd852917899;
array[11901]=30'd852917899;
array[11902]=30'd852917899;
array[11903]=30'd852917899;
array[11904]=30'd852917899;
array[11905]=30'd852917899;
array[11906]=30'd852917899;
array[11907]=30'd873911932;
array[11908]=30'd873911932;
array[11909]=30'd873911932;
array[11910]=30'd873911932;
array[11911]=30'd873911932;
array[11912]=30'd873911932;
array[11913]=30'd873911932;
array[11914]=30'd900139626;
array[11915]=30'd898098744;
array[11916]=30'd875034136;
array[11917]=30'd764964292;
array[11918]=30'd794289609;
array[11919]=30'd794289609;
array[11920]=30'd794289609;
array[11921]=30'd820487650;
array[11922]=30'd820487650;
array[11923]=30'd844591615;
array[11924]=30'd862402083;
array[11925]=30'd867617357;
array[11926]=30'd852917899;
array[11927]=30'd873911932;
array[11928]=30'd873911932;
array[11929]=30'd873911932;
array[11930]=30'd873911932;
array[11931]=30'd873911932;
array[11932]=30'd873911932;
array[11933]=30'd873911932;
array[11934]=30'd873911932;
array[11935]=30'd873911932;
array[11936]=30'd852917899;
array[11937]=30'd873911932;
array[11938]=30'd873911932;
array[11939]=30'd873911932;
array[11940]=30'd852917899;
array[11941]=30'd852917899;
array[11942]=30'd852917899;
array[11943]=30'd852917899;
array[11944]=30'd581297788;
array[11945]=30'd636841618;
array[11946]=30'd644165300;
array[11947]=30'd485848753;
array[11948]=30'd653646508;
array[11949]=30'd625391195;
array[11950]=30'd941029952;
array[11951]=30'd757545539;
array[11952]=30'd757545539;
array[11953]=30'd721911330;
array[11954]=30'd472349226;
array[11955]=30'd352820791;
array[11956]=30'd595020337;
array[11957]=30'd916923947;
array[11958]=30'd959928886;
array[11959]=30'd985089582;
array[11960]=30'd985089582;
array[11961]=30'd959928886;
array[11962]=30'd959928886;
array[11963]=30'd959928886;
array[11964]=30'd941029952;
array[11965]=30'd757545539;
array[11966]=30'd809995819;
array[11967]=30'd721911330;
array[11968]=30'd679964212;
array[11969]=30'd721911330;
array[11970]=30'd679964212;
array[11971]=30'd721911330;
array[11972]=30'd916923947;
array[11973]=30'd959928886;
array[11974]=30'd959928886;
array[11975]=30'd935829023;
array[11976]=30'd721911330;
array[11977]=30'd511088198;
array[11978]=30'd626373227;
array[11979]=30'd452327079;
array[11980]=30'd644165300;
array[11981]=30'd632612564;
array[11982]=30'd596983478;
array[11983]=30'd557159098;
array[11984]=30'd632612564;
array[11985]=30'd549823127;
array[11986]=30'd852917899;
array[11987]=30'd852917899;
array[11988]=30'd852917899;
array[11989]=30'd852917899;
array[11990]=30'd852917899;
array[11991]=30'd852917899;
array[11992]=30'd852917899;
array[11993]=30'd852917899;
array[11994]=30'd852917899;
array[11995]=30'd852917899;
array[11996]=30'd852917899;
array[11997]=30'd852917899;
array[11998]=30'd852917899;
array[11999]=30'd852917899;
array[12000]=30'd852917899;
array[12001]=30'd873911932;
array[12002]=30'd852917899;
array[12003]=30'd873911932;
array[12004]=30'd873911932;
array[12005]=30'd873911932;
array[12006]=30'd873911932;
array[12007]=30'd873911932;
array[12008]=30'd873911932;
array[12009]=30'd873911932;
array[12010]=30'd900139626;
array[12011]=30'd959928886;
array[12012]=30'd926429685;
array[12013]=30'd820487650;
array[12014]=30'd844591615;
array[12015]=30'd910663171;
array[12016]=30'd844591615;
array[12017]=30'd862402083;
array[12018]=30'd862402083;
array[12019]=30'd887567935;
array[12020]=30'd867617357;
array[12021]=30'd873911932;
array[12022]=30'd873911932;
array[12023]=30'd873911932;
array[12024]=30'd873911932;
array[12025]=30'd873911932;
array[12026]=30'd873911932;
array[12027]=30'd873911932;
array[12028]=30'd873911932;
array[12029]=30'd873911932;
array[12030]=30'd873911932;
array[12031]=30'd873911932;
array[12032]=30'd873911932;
array[12033]=30'd873911932;
array[12034]=30'd873911932;
array[12035]=30'd873911932;
array[12036]=30'd873911932;
array[12037]=30'd873911932;
array[12038]=30'd852917899;
array[12039]=30'd852917899;
array[12040]=30'd593947240;
array[12041]=30'd636841618;
array[12042]=30'd644165300;
array[12043]=30'd485848753;
array[12044]=30'd653646508;
array[12045]=30'd560346760;
array[12046]=30'd840392271;
array[12047]=30'd809995819;
array[12048]=30'd501707283;
array[12049]=30'd395804188;
array[12050]=30'd721911330;
array[12051]=30'd778555959;
array[12052]=30'd556237353;
array[12053]=30'd472349226;
array[12054]=30'd941029952;
array[12055]=30'd985089582;
array[12056]=30'd959928886;
array[12057]=30'd959928886;
array[12058]=30'd959928886;
array[12059]=30'd959928886;
array[12060]=30'd959928886;
array[12061]=30'd642228804;
array[12062]=30'd352820791;
array[12063]=30'd617068069;
array[12064]=30'd679964212;
array[12065]=30'd472349226;
array[12066]=30'd252147238;
array[12067]=30'd501707283;
array[12068]=30'd679964212;
array[12069]=30'd887567935;
array[12070]=30'd959928886;
array[12071]=30'd916923947;
array[12072]=30'd794232376;
array[12073]=30'd581297788;
array[12074]=30'd636841618;
array[12075]=30'd452327079;
array[12076]=30'd644165300;
array[12077]=30'd644165300;
array[12078]=30'd596983478;
array[12079]=30'd557159098;
array[12080]=30'd644165300;
array[12081]=30'd549823127;
array[12082]=30'd873911932;
array[12083]=30'd852917899;
array[12084]=30'd852917899;
array[12085]=30'd873911932;
array[12086]=30'd852917899;
array[12087]=30'd873911932;
array[12088]=30'd873911932;
array[12089]=30'd873911932;
array[12090]=30'd873911932;
array[12091]=30'd852917899;
array[12092]=30'd852917899;
array[12093]=30'd852917899;
array[12094]=30'd852917899;
array[12095]=30'd852917899;
array[12096]=30'd852917899;
array[12097]=30'd873911932;
array[12098]=30'd873911932;
array[12099]=30'd873911932;
array[12100]=30'd873911932;
array[12101]=30'd873911932;
array[12102]=30'd873911932;
array[12103]=30'd873911932;
array[12104]=30'd873911932;
array[12105]=30'd900139626;
array[12106]=30'd921150041;
array[12107]=30'd1004004888;
array[12108]=30'd855119352;
array[12109]=30'd778567150;
array[12110]=30'd935829023;
array[12111]=30'd967280137;
array[12112]=30'd855119352;
array[12113]=30'd862402083;
array[12114]=30'd916923947;
array[12115]=30'd935829023;
array[12116]=30'd862402083;
array[12117]=30'd887567935;
array[12118]=30'd867617357;
array[12119]=30'd873911932;
array[12120]=30'd873911932;
array[12121]=30'd873911932;
array[12122]=30'd873911932;
array[12123]=30'd873911932;
array[12124]=30'd873911932;
array[12125]=30'd873911932;
array[12126]=30'd873911932;
array[12127]=30'd873911932;
array[12128]=30'd873911932;
array[12129]=30'd873911932;
array[12130]=30'd873911932;
array[12131]=30'd873911932;
array[12132]=30'd873911932;
array[12133]=30'd873911932;
array[12134]=30'd852917899;
array[12135]=30'd852917899;
array[12136]=30'd625391195;
array[12137]=30'd636841618;
array[12138]=30'd644165300;
array[12139]=30'd444947126;
array[12140]=30'd653646508;
array[12141]=30'd604360306;
array[12142]=30'd840392271;
array[12143]=30'd352820791;
array[12144]=30'd617068069;
array[12145]=30'd935829023;
array[12146]=30'd959928886;
array[12147]=30'd959928886;
array[12148]=30'd959928886;
array[12149]=30'd887567935;
array[12150]=30'd959928886;
array[12151]=30'd959928886;
array[12152]=30'd959928886;
array[12153]=30'd959928886;
array[12154]=30'd959928886;
array[12155]=30'd959928886;
array[12156]=30'd959928886;
array[12157]=30'd862402083;
array[12158]=30'd916923947;
array[12159]=30'd959928886;
array[12160]=30'd959928886;
array[12161]=30'd959928886;
array[12162]=30'd809995819;
array[12163]=30'd395804188;
array[12164]=30'd308796939;
array[12165]=30'd809995819;
array[12166]=30'd959928886;
array[12167]=30'd941029952;
array[12168]=30'd757545539;
array[12169]=30'd604360306;
array[12170]=30'd636841618;
array[12171]=30'd461756049;
array[12172]=30'd515208870;
array[12173]=30'd644165300;
array[12174]=30'd557159098;
array[12175]=30'd596983478;
array[12176]=30'd644165300;
array[12177]=30'd653676161;
array[12178]=30'd887567935;
array[12179]=30'd867617357;
array[12180]=30'd900139626;
array[12181]=30'd900139626;
array[12182]=30'd941029952;
array[12183]=30'd941029952;
array[12184]=30'd941029952;
array[12185]=30'd941029952;
array[12186]=30'd900139626;
array[12187]=30'd873911932;
array[12188]=30'd873911932;
array[12189]=30'd873911932;
array[12190]=30'd852917899;
array[12191]=30'd852917899;
array[12192]=30'd852917899;
array[12193]=30'd852917899;
array[12194]=30'd873911932;
array[12195]=30'd873911932;
array[12196]=30'd873911932;
array[12197]=30'd873911932;
array[12198]=30'd873911932;
array[12199]=30'd873911932;
array[12200]=30'd873911932;
array[12201]=30'd900139626;
array[12202]=30'd959928886;
array[12203]=30'd926429685;
array[12204]=30'd785935846;
array[12205]=30'd844591615;
array[12206]=30'd967280137;
array[12207]=30'd950544914;
array[12208]=30'd752351692;
array[12209]=30'd820487650;
array[12210]=30'd935829023;
array[12211]=30'd926429685;
array[12212]=30'd752351692;
array[12213]=30'd844591615;
array[12214]=30'd862402083;
array[12215]=30'd873911932;
array[12216]=30'd873911932;
array[12217]=30'd873911932;
array[12218]=30'd873911932;
array[12219]=30'd873911932;
array[12220]=30'd873911932;
array[12221]=30'd873911932;
array[12222]=30'd873911932;
array[12223]=30'd873911932;
array[12224]=30'd873911932;
array[12225]=30'd873911932;
array[12226]=30'd873911932;
array[12227]=30'd873911932;
array[12228]=30'd873911932;
array[12229]=30'd873911932;
array[12230]=30'd873911932;
array[12231]=30'd873911932;
array[12232]=30'd684081775;
array[12233]=30'd609598119;
array[12234]=30'd644165300;
array[12235]=30'd485848753;
array[12236]=30'd653646508;
array[12237]=30'd560346760;
array[12238]=30'd642228804;
array[12239]=30'd617068069;
array[12240]=30'd959928886;
array[12241]=30'd959928886;
array[12242]=30'd959928886;
array[12243]=30'd959928886;
array[12244]=30'd959928886;
array[12245]=30'd985089582;
array[12246]=30'd959928886;
array[12247]=30'd959928886;
array[12248]=30'd959928886;
array[12249]=30'd959928886;
array[12250]=30'd959928886;
array[12251]=30'd959928886;
array[12252]=30'd959928886;
array[12253]=30'd959928886;
array[12254]=30'd959928886;
array[12255]=30'd959928886;
array[12256]=30'd959928886;
array[12257]=30'd959928886;
array[12258]=30'd959928886;
array[12259]=30'd916923947;
array[12260]=30'd556237353;
array[12261]=30'd395804188;
array[12262]=30'd959928886;
array[12263]=30'd941029952;
array[12264]=30'd666281541;
array[12265]=30'd626373227;
array[12266]=30'd609598119;
array[12267]=30'd397801110;
array[12268]=30'd557159098;
array[12269]=30'd644165300;
array[12270]=30'd515208870;
array[12271]=30'd596983478;
array[12272]=30'd609598119;
array[12273]=30'd709314133;
array[12274]=30'd941029952;
array[12275]=30'd916923947;
array[12276]=30'd910663171;
array[12277]=30'd875034136;
array[12278]=30'd888658404;
array[12279]=30'd888658404;
array[12280]=30'd904416730;
array[12281]=30'd946320871;
array[12282]=30'd967280137;
array[12283]=30'd941029952;
array[12284]=30'd873911932;
array[12285]=30'd873911932;
array[12286]=30'd852917899;
array[12287]=30'd873911932;
array[12288]=30'd873911932;
array[12289]=30'd873911932;
array[12290]=30'd873911932;
array[12291]=30'd873911932;
array[12292]=30'd873911932;
array[12293]=30'd873911932;
array[12294]=30'd873911932;
array[12295]=30'd873911932;
array[12296]=30'd873911932;
array[12297]=30'd900139626;
array[12298]=30'd935829023;
array[12299]=30'd785935846;
array[12300]=30'd785935846;
array[12301]=30'd890710541;
array[12302]=30'd935829023;
array[12303]=30'd926429685;
array[12304]=30'd764964292;
array[12305]=30'd794289609;
array[12306]=30'd910663171;
array[12307]=30'd987238908;
array[12308]=30'd764964292;
array[12309]=30'd794289609;
array[12310]=30'd890710541;
array[12311]=30'd867617357;
array[12312]=30'd873911932;
array[12313]=30'd873911932;
array[12314]=30'd873911932;
array[12315]=30'd873911932;
array[12316]=30'd873911932;
array[12317]=30'd873911932;
array[12318]=30'd873911932;
array[12319]=30'd873911932;
array[12320]=30'd873911932;
array[12321]=30'd873911932;
array[12322]=30'd873911932;
array[12323]=30'd873911932;
array[12324]=30'd873911932;
array[12325]=30'd873911932;
array[12326]=30'd873911932;
array[12327]=30'd873911932;
array[12328]=30'd709304966;
array[12329]=30'd609598119;
array[12330]=30'd644165300;
array[12331]=30'd485848753;
array[12332]=30'd653646508;
array[12333]=30'd560346760;
array[12334]=30'd941029952;
array[12335]=30'd941029952;
array[12336]=30'd959928886;
array[12337]=30'd959928886;
array[12338]=30'd959928886;
array[12339]=30'd959928886;
array[12340]=30'd959928886;
array[12341]=30'd959928886;
array[12342]=30'd959928886;
array[12343]=30'd959928886;
array[12344]=30'd959928886;
array[12345]=30'd959928886;
array[12346]=30'd959928886;
array[12347]=30'd959928886;
array[12348]=30'd959928886;
array[12349]=30'd959928886;
array[12350]=30'd959928886;
array[12351]=30'd959928886;
array[12352]=30'd959928886;
array[12353]=30'd959928886;
array[12354]=30'd959928886;
array[12355]=30'd959928886;
array[12356]=30'd941029952;
array[12357]=30'd809995819;
array[12358]=30'd959928886;
array[12359]=30'd941029952;
array[12360]=30'd593947240;
array[12361]=30'd636841618;
array[12362]=30'd609598119;
array[12363]=30'd397801110;
array[12364]=30'd596983478;
array[12365]=30'd644165300;
array[12366]=30'd515208870;
array[12367]=30'd644165300;
array[12368]=30'd557159098;
array[12369]=30'd757545539;
array[12370]=30'd875034136;
array[12371]=30'd785935846;
array[12372]=30'd764964292;
array[12373]=30'd764964292;
array[12374]=30'd764964292;
array[12375]=30'd782796193;
array[12376]=30'd782796193;
array[12377]=30'd782796193;
array[12378]=30'd929554891;
array[12379]=30'd967280137;
array[12380]=30'd887567935;
array[12381]=30'd873911932;
array[12382]=30'd873911932;
array[12383]=30'd852917899;
array[12384]=30'd873911932;
array[12385]=30'd873911932;
array[12386]=30'd873911932;
array[12387]=30'd873911932;
array[12388]=30'd873911932;
array[12389]=30'd873911932;
array[12390]=30'd873911932;
array[12391]=30'd873911932;
array[12392]=30'd873911932;
array[12393]=30'd900139626;
array[12394]=30'd857219651;
array[12395]=30'd809995819;
array[12396]=30'd862402083;
array[12397]=30'd887567935;
array[12398]=30'd935829023;
array[12399]=30'd926429685;
array[12400]=30'd752351692;
array[12401]=30'd820487650;
array[12402]=30'd890710541;
array[12403]=30'd950544914;
array[12404]=30'd785935846;
array[12405]=30'd820487650;
array[12406]=30'd862402083;
array[12407]=30'd867617357;
array[12408]=30'd873911932;
array[12409]=30'd900139626;
array[12410]=30'd873911932;
array[12411]=30'd873911932;
array[12412]=30'd873911932;
array[12413]=30'd873911932;
array[12414]=30'd873911932;
array[12415]=30'd873911932;
array[12416]=30'd873911932;
array[12417]=30'd873911932;
array[12418]=30'd873911932;
array[12419]=30'd873911932;
array[12420]=30'd873911932;
array[12421]=30'd873911932;
array[12422]=30'd873911932;
array[12423]=30'd873911932;
array[12424]=30'd773214847;
array[12425]=30'd549823127;
array[12426]=30'd644165300;
array[12427]=30'd444947126;
array[12428]=30'd653646508;
array[12429]=30'd527847013;
array[12430]=30'd840392271;
array[12431]=30'd887567935;
array[12432]=30'd887567935;
array[12433]=30'd916923947;
array[12434]=30'd941029952;
array[12435]=30'd916923947;
array[12436]=30'd959928886;
array[12437]=30'd959928886;
array[12438]=30'd959928886;
array[12439]=30'd959928886;
array[12440]=30'd959928886;
array[12441]=30'd959928886;
array[12442]=30'd959928886;
array[12443]=30'd959928886;
array[12444]=30'd959928886;
array[12445]=30'd959928886;
array[12446]=30'd959928886;
array[12447]=30'd959928886;
array[12448]=30'd959928886;
array[12449]=30'd887567935;
array[12450]=30'd959928886;
array[12451]=30'd941029952;
array[12452]=30'd887567935;
array[12453]=30'd959928886;
array[12454]=30'd941029952;
array[12455]=30'd887567935;
array[12456]=30'd553016910;
array[12457]=30'd636841618;
array[12458]=30'd557159098;
array[12459]=30'd427157133;
array[12460]=30'd644165300;
array[12461]=30'd644165300;
array[12462]=30'd515208870;
array[12463]=30'd644165300;
array[12464]=30'd522581659;
array[12465]=30'd804758111;
array[12466]=30'd832058842;
array[12467]=30'd785935846;
array[12468]=30'd811098555;
array[12469]=30'd832058842;
array[12470]=30'd869807552;
array[12471]=30'd906527146;
array[12472]=30'd906527146;
array[12473]=30'd833137031;
array[12474]=30'd782796193;
array[12475]=30'd946320871;
array[12476]=30'd935829023;
array[12477]=30'd867617357;
array[12478]=30'd873911932;
array[12479]=30'd852917899;
array[12480]=30'd873911932;
array[12481]=30'd873911932;
array[12482]=30'd873911932;
array[12483]=30'd873911932;
array[12484]=30'd873911932;
array[12485]=30'd873911932;
array[12486]=30'd873911932;
array[12487]=30'd873911932;
array[12488]=30'd900139626;
array[12489]=30'd900139626;
array[12490]=30'd900139626;
array[12491]=30'd887567935;
array[12492]=30'd867617357;
array[12493]=30'd900139626;
array[12494]=30'd921150041;
array[12495]=30'd857219651;
array[12496]=30'd778567150;
array[12497]=30'd870795757;
array[12498]=30'd887567935;
array[12499]=30'd887567935;
array[12500]=30'd887567935;
array[12501]=30'd862402083;
array[12502]=30'd867617357;
array[12503]=30'd873911932;
array[12504]=30'd873911932;
array[12505]=30'd873911932;
array[12506]=30'd873911932;
array[12507]=30'd873911932;
array[12508]=30'd873911932;
array[12509]=30'd873911932;
array[12510]=30'd873911932;
array[12511]=30'd873911932;
array[12512]=30'd873911932;
array[12513]=30'd873911932;
array[12514]=30'd873911932;
array[12515]=30'd873911932;
array[12516]=30'd873911932;
array[12517]=30'd873911932;
array[12518]=30'd873911932;
array[12519]=30'd873911932;
array[12520]=30'd815162003;
array[12521]=30'd522581659;
array[12522]=30'd644165300;
array[12523]=30'd452327079;
array[12524]=30'd653646508;
array[12525]=30'd625391195;
array[12526]=30'd941029952;
array[12527]=30'd959928886;
array[12528]=30'd887567935;
array[12529]=30'd959928886;
array[12530]=30'd959928886;
array[12531]=30'd959928886;
array[12532]=30'd959928886;
array[12533]=30'd959928886;
array[12534]=30'd959928886;
array[12535]=30'd959928886;
array[12536]=30'd959928886;
array[12537]=30'd959928886;
array[12538]=30'd959928886;
array[12539]=30'd959928886;
array[12540]=30'd959928886;
array[12541]=30'd959928886;
array[12542]=30'd959928886;
array[12543]=30'd959928886;
array[12544]=30'd916923947;
array[12545]=30'd941029952;
array[12546]=30'd959928886;
array[12547]=30'd887567935;
array[12548]=30'd959928886;
array[12549]=30'd959928886;
array[12550]=30'd840392271;
array[12551]=30'd862402083;
array[12552]=30'd527847013;
array[12553]=30'd636841618;
array[12554]=30'd515208870;
array[12555]=30'd496374434;
array[12556]=30'd644165300;
array[12557]=30'd596983478;
array[12558]=30'd557159098;
array[12559]=30'd644165300;
array[12560]=30'd560346760;
array[12561]=30'd857219651;
array[12562]=30'd785935846;
array[12563]=30'd869807552;
array[12564]=30'd888658404;
array[12565]=30'd855119352;
array[12566]=30'd869807552;
array[12567]=30'd811098555;
array[12568]=30'd782796193;
array[12569]=30'd849905057;
array[12570]=30'd833137031;
array[12571]=30'd869807552;
array[12572]=30'd967280137;
array[12573]=30'd887567935;
array[12574]=30'd867617357;
array[12575]=30'd852917899;
array[12576]=30'd873911932;
array[12577]=30'd873911932;
array[12578]=30'd873911932;
array[12579]=30'd873911932;
array[12580]=30'd873911932;
array[12581]=30'd873911932;
array[12582]=30'd873911932;
array[12583]=30'd900139626;
array[12584]=30'd873911932;
array[12585]=30'd873911932;
array[12586]=30'd873911932;
array[12587]=30'd873911932;
array[12588]=30'd873911932;
array[12589]=30'd873911932;
array[12590]=30'd900139626;
array[12591]=30'd900139626;
array[12592]=30'd887567935;
array[12593]=30'd887567935;
array[12594]=30'd900139626;
array[12595]=30'd873911932;
array[12596]=30'd900139626;
array[12597]=30'd873911932;
array[12598]=30'd873911932;
array[12599]=30'd873911932;
array[12600]=30'd873911932;
array[12601]=30'd873911932;
array[12602]=30'd873911932;
array[12603]=30'd873911932;
array[12604]=30'd873911932;
array[12605]=30'd873911932;
array[12606]=30'd873911932;
array[12607]=30'd873911932;
array[12608]=30'd873911932;
array[12609]=30'd873911932;
array[12610]=30'd873911932;
array[12611]=30'd873911932;
array[12612]=30'd873911932;
array[12613]=30'd873911932;
array[12614]=30'd873911932;
array[12615]=30'd873911932;
array[12616]=30'd852917899;
array[12617]=30'd522581659;
array[12618]=30'd636841618;
array[12619]=30'd452327079;
array[12620]=30'd609598119;
array[12621]=30'd740735615;
array[12622]=30'd959928886;
array[12623]=30'd959928886;
array[12624]=30'd959928886;
array[12625]=30'd959928886;
array[12626]=30'd959928886;
array[12627]=30'd959928886;
array[12628]=30'd959928886;
array[12629]=30'd959928886;
array[12630]=30'd959928886;
array[12631]=30'd959928886;
array[12632]=30'd959928886;
array[12633]=30'd959928886;
array[12634]=30'd959928886;
array[12635]=30'd959928886;
array[12636]=30'd959928886;
array[12637]=30'd959928886;
array[12638]=30'd959928886;
array[12639]=30'd959928886;
array[12640]=30'd959928886;
array[12641]=30'd959928886;
array[12642]=30'd959928886;
array[12643]=30'd959928886;
array[12644]=30'd959928886;
array[12645]=30'd959928886;
array[12646]=30'd941029952;
array[12647]=30'd794232376;
array[12648]=30'd581297788;
array[12649]=30'd636841618;
array[12650]=30'd461756049;
array[12651]=30'd557159098;
array[12652]=30'd644165300;
array[12653]=30'd515208870;
array[12654]=30'd609598119;
array[12655]=30'd609598119;
array[12656]=30'd653676161;
array[12657]=30'd820526616;
array[12658]=30'd785935846;
array[12659]=30'd904416730;
array[12660]=30'd855119352;
array[12661]=30'd778567150;
array[12662]=30'd764964292;
array[12663]=30'd782796193;
array[12664]=30'd782796193;
array[12665]=30'd768126344;
array[12666]=30'd833137031;
array[12667]=30'd782796193;
array[12668]=30'd929554891;
array[12669]=30'd910663171;
array[12670]=30'd867617357;
array[12671]=30'd873911932;
array[12672]=30'd900139626;
array[12673]=30'd900139626;
array[12674]=30'd900139626;
array[12675]=30'd873911932;
array[12676]=30'd873911932;
array[12677]=30'd900139626;
array[12678]=30'd873911932;
array[12679]=30'd873911932;
array[12680]=30'd900139626;
array[12681]=30'd873911932;
array[12682]=30'd900139626;
array[12683]=30'd873911932;
array[12684]=30'd873911932;
array[12685]=30'd900139626;
array[12686]=30'd900139626;
array[12687]=30'd873911932;
array[12688]=30'd873911932;
array[12689]=30'd873911932;
array[12690]=30'd873911932;
array[12691]=30'd873911932;
array[12692]=30'd873911932;
array[12693]=30'd873911932;
array[12694]=30'd873911932;
array[12695]=30'd873911932;
array[12696]=30'd873911932;
array[12697]=30'd873911932;
array[12698]=30'd873911932;
array[12699]=30'd873911932;
array[12700]=30'd873911932;
array[12701]=30'd873911932;
array[12702]=30'd873911932;
array[12703]=30'd873911932;
array[12704]=30'd873911932;
array[12705]=30'd873911932;
array[12706]=30'd873911932;
array[12707]=30'd873911932;
array[12708]=30'd873911932;
array[12709]=30'd873911932;
array[12710]=30'd873911932;
array[12711]=30'd873911932;
array[12712]=30'd852917899;
array[12713]=30'd604360306;
array[12714]=30'd636841618;
array[12715]=30'd461756049;
array[12716]=30'd557159098;
array[12717]=30'd821480030;
array[12718]=30'd959928886;
array[12719]=30'd959928886;
array[12720]=30'd959928886;
array[12721]=30'd959928886;
array[12722]=30'd959928886;
array[12723]=30'd959928886;
array[12724]=30'd959928886;
array[12725]=30'd959928886;
array[12726]=30'd959928886;
array[12727]=30'd959928886;
array[12728]=30'd959928886;
array[12729]=30'd959928886;
array[12730]=30'd959928886;
array[12731]=30'd959928886;
array[12732]=30'd959928886;
array[12733]=30'd959928886;
array[12734]=30'd959928886;
array[12735]=30'd985089582;
array[12736]=30'd959928886;
array[12737]=30'd959928886;
array[12738]=30'd959928886;
array[12739]=30'd959928886;
array[12740]=30'd959928886;
array[12741]=30'd959928886;
array[12742]=30'd941029952;
array[12743]=30'd740728401;
array[12744]=30'd626373227;
array[12745]=30'd609598119;
array[12746]=30'd427157133;
array[12747]=30'd609598119;
array[12748]=30'd644165300;
array[12749]=30'd461756049;
array[12750]=30'd653646508;
array[12751]=30'd557159098;
array[12752]=30'd709304966;
array[12753]=30'd820526616;
array[12754]=30'd832058842;
array[12755]=30'd888658404;
array[12756]=30'd855119352;
array[12757]=30'd785935846;
array[12758]=30'd869807552;
array[12759]=30'd945318330;
array[12760]=30'd849905057;
array[12761]=30'd782796193;
array[12762]=30'd885566856;
array[12763]=30'd782796193;
array[12764]=30'd869807552;
array[12765]=30'd946320871;
array[12766]=30'd867617357;
array[12767]=30'd873911932;
array[12768]=30'd887567935;
array[12769]=30'd916923947;
array[12770]=30'd887567935;
array[12771]=30'd887567935;
array[12772]=30'd900139626;
array[12773]=30'd900139626;
array[12774]=30'd873911932;
array[12775]=30'd873911932;
array[12776]=30'd900139626;
array[12777]=30'd900139626;
array[12778]=30'd900139626;
array[12779]=30'd900139626;
array[12780]=30'd873911932;
array[12781]=30'd873911932;
array[12782]=30'd900139626;
array[12783]=30'd873911932;
array[12784]=30'd873911932;
array[12785]=30'd873911932;
array[12786]=30'd900139626;
array[12787]=30'd900139626;
array[12788]=30'd873911932;
array[12789]=30'd873911932;
array[12790]=30'd873911932;
array[12791]=30'd873911932;
array[12792]=30'd873911932;
array[12793]=30'd873911932;
array[12794]=30'd873911932;
array[12795]=30'd900139626;
array[12796]=30'd873911932;
array[12797]=30'd900139626;
array[12798]=30'd873911932;
array[12799]=30'd873911932;
array[12800]=30'd873911932;
array[12801]=30'd873911932;
array[12802]=30'd873911932;
array[12803]=30'd873911932;
array[12804]=30'd873911932;
array[12805]=30'd873911932;
array[12806]=30'd873911932;
array[12807]=30'd873911932;
array[12808]=30'd873911932;
array[12809]=30'd710295175;
array[12810]=30'd581297788;
array[12811]=30'd461756049;
array[12812]=30'd609598119;
array[12813]=30'd821480030;
array[12814]=30'd959928886;
array[12815]=30'd959928886;
array[12816]=30'd959928886;
array[12817]=30'd959928886;
array[12818]=30'd959928886;
array[12819]=30'd959928886;
array[12820]=30'd941029952;
array[12821]=30'd862402083;
array[12822]=30'd916923947;
array[12823]=30'd941029952;
array[12824]=30'd959928886;
array[12825]=30'd959928886;
array[12826]=30'd959928886;
array[12827]=30'd959928886;
array[12828]=30'd959928886;
array[12829]=30'd916923947;
array[12830]=30'd862402083;
array[12831]=30'd959928886;
array[12832]=30'd959928886;
array[12833]=30'd959928886;
array[12834]=30'd959928886;
array[12835]=30'd959928886;
array[12836]=30'd959928886;
array[12837]=30'd941029952;
array[12838]=30'd941029952;
array[12839]=30'd625391195;
array[12840]=30'd636841618;
array[12841]=30'd609598119;
array[12842]=30'd496374434;
array[12843]=30'd636841618;
array[12844]=30'd549823127;
array[12845]=30'd461756049;
array[12846]=30'd636841618;
array[12847]=30'd522581659;
array[12848]=30'd783791725;
array[12849]=30'd778567150;
array[12850]=30'd869807552;
array[12851]=30'd910663171;
array[12852]=30'd875034136;
array[12853]=30'd785935846;
array[12854]=30'd849905057;
array[12855]=30'd945318330;
array[12856]=30'd869807552;
array[12857]=30'd782796193;
array[12858]=30'd849905057;
array[12859]=30'd833137031;
array[12860]=30'd811098555;
array[12861]=30'd946320871;
array[12862]=30'd887567935;
array[12863]=30'd873911932;
array[12864]=30'd862402083;
array[12865]=30'd875034136;
array[12866]=30'd844591615;
array[12867]=30'd890710541;
array[12868]=30'd887567935;
array[12869]=30'd900139626;
array[12870]=30'd900139626;
array[12871]=30'd873911932;
array[12872]=30'd873911932;
array[12873]=30'd873911932;
array[12874]=30'd873911932;
array[12875]=30'd900139626;
array[12876]=30'd873911932;
array[12877]=30'd873911932;
array[12878]=30'd900139626;
array[12879]=30'd900139626;
array[12880]=30'd900139626;
array[12881]=30'd873911932;
array[12882]=30'd873911932;
array[12883]=30'd873911932;
array[12884]=30'd873911932;
array[12885]=30'd873911932;
array[12886]=30'd900139626;
array[12887]=30'd900139626;
array[12888]=30'd900139626;
array[12889]=30'd900139626;
array[12890]=30'd900139626;
array[12891]=30'd900139626;
array[12892]=30'd873911932;
array[12893]=30'd900139626;
array[12894]=30'd900139626;
array[12895]=30'd873911932;
array[12896]=30'd873911932;
array[12897]=30'd873911932;
array[12898]=30'd873911932;
array[12899]=30'd900139626;
array[12900]=30'd900139626;
array[12901]=30'd873911932;
array[12902]=30'd873911932;
array[12903]=30'd873911932;
array[12904]=30'd873911932;
array[12905]=30'd792127082;
array[12906]=30'd527847013;
array[12907]=30'd461756049;
array[12908]=30'd653646508;
array[12909]=30'd684081775;
array[12910]=30'd959928886;
array[12911]=30'd959928886;
array[12912]=30'd959928886;
array[12913]=30'd959928886;
array[12914]=30'd959928886;
array[12915]=30'd959928886;
array[12916]=30'd959928886;
array[12917]=30'd916923947;
array[12918]=30'd862402083;
array[12919]=30'd794232376;
array[12920]=30'd794232376;
array[12921]=30'd794232376;
array[12922]=30'd809995819;
array[12923]=30'd794232376;
array[12924]=30'd757545539;
array[12925]=30'd809995819;
array[12926]=30'd916923947;
array[12927]=30'd959928886;
array[12928]=30'd959928886;
array[12929]=30'd959928886;
array[12930]=30'd959928886;
array[12931]=30'd959928886;
array[12932]=30'd959928886;
array[12933]=30'd941029952;
array[12934]=30'd916923947;
array[12935]=30'd553016910;
array[12936]=30'd666201723;
array[12937]=30'd549823127;
array[12938]=30'd609598119;
array[12939]=30'd609598119;
array[12940]=30'd427157133;
array[12941]=30'd522581659;
array[12942]=30'd653646508;
array[12943]=30'd522581659;
array[12944]=30'd840392271;
array[12945]=30'd778567150;
array[12946]=30'd869807552;
array[12947]=30'd910663171;
array[12948]=30'd875034136;
array[12949]=30'd785935846;
array[12950]=30'd811098555;
array[12951]=30'd906527146;
array[12952]=30'd811098555;
array[12953]=30'd764964292;
array[12954]=30'd849905057;
array[12955]=30'd833137031;
array[12956]=30'd811098555;
array[12957]=30'd888658404;
array[12958]=30'd887567935;
array[12959]=30'd873911932;
array[12960]=30'd910663171;
array[12961]=30'd888658404;
array[12962]=30'd832058842;
array[12963]=30'd890710541;
array[12964]=30'd887567935;
array[12965]=30'd900139626;
array[12966]=30'd873911932;
array[12967]=30'd873911932;
array[12968]=30'd900139626;
array[12969]=30'd900139626;
array[12970]=30'd900139626;
array[12971]=30'd900139626;
array[12972]=30'd900139626;
array[12973]=30'd873911932;
array[12974]=30'd900139626;
array[12975]=30'd900139626;
array[12976]=30'd900139626;
array[12977]=30'd873911932;
array[12978]=30'd900139626;
array[12979]=30'd900139626;
array[12980]=30'd900139626;
array[12981]=30'd900139626;
array[12982]=30'd900139626;
array[12983]=30'd900139626;
array[12984]=30'd900139626;
array[12985]=30'd900139626;
array[12986]=30'd900139626;
array[12987]=30'd873911932;
array[12988]=30'd900139626;
array[12989]=30'd900139626;
array[12990]=30'd900139626;
array[12991]=30'd873911932;
array[12992]=30'd900139626;
array[12993]=30'd900139626;
array[12994]=30'd900139626;
array[12995]=30'd900139626;
array[12996]=30'd900139626;
array[12997]=30'd900139626;
array[12998]=30'd873911932;
array[12999]=30'd873911932;
array[13000]=30'd873911932;
array[13001]=30'd852917899;
array[13002]=30'd503733877;
array[13003]=30'd486913656;
array[13004]=30'd674612899;
array[13005]=30'd604360306;
array[13006]=30'd804758111;
array[13007]=30'd959928886;
array[13008]=30'd959928886;
array[13009]=30'd959928886;
array[13010]=30'd959928886;
array[13011]=30'd959928886;
array[13012]=30'd959928886;
array[13013]=30'd959928886;
array[13014]=30'd959928886;
array[13015]=30'd959928886;
array[13016]=30'd985089582;
array[13017]=30'd985089582;
array[13018]=30'd959928886;
array[13019]=30'd959928886;
array[13020]=30'd959928886;
array[13021]=30'd959928886;
array[13022]=30'd959928886;
array[13023]=30'd959928886;
array[13024]=30'd959928886;
array[13025]=30'd985089582;
array[13026]=30'd959928886;
array[13027]=30'd959928886;
array[13028]=30'd959928886;
array[13029]=30'd941029952;
array[13030]=30'd867617357;
array[13031]=30'd527847013;
array[13032]=30'd636841618;
array[13033]=30'd444947126;
array[13034]=30'd644165300;
array[13035]=30'd557159098;
array[13036]=30'd364251806;
array[13037]=30'd557159098;
array[13038]=30'd636841618;
array[13039]=30'd593947240;
array[13040]=30'd887567935;
array[13041]=30'd785935846;
array[13042]=30'd869807552;
array[13043]=30'd967280137;
array[13044]=30'd875034136;
array[13045]=30'd785935846;
array[13046]=30'd811098555;
array[13047]=30'd945318330;
array[13048]=30'd869807552;
array[13049]=30'd811098555;
array[13050]=30'd849905057;
array[13051]=30'd782796193;
array[13052]=30'd832058842;
array[13053]=30'd910663171;
array[13054]=30'd867617357;
array[13055]=30'd873911932;
array[13056]=30'd875034136;
array[13057]=30'd855119352;
array[13058]=30'd832058842;
array[13059]=30'd870795757;
array[13060]=30'd887567935;
array[13061]=30'd887567935;
array[13062]=30'd900139626;
array[13063]=30'd900139626;
array[13064]=30'd900139626;
array[13065]=30'd900139626;
array[13066]=30'd900139626;
array[13067]=30'd900139626;
array[13068]=30'd900139626;
array[13069]=30'd900139626;
array[13070]=30'd900139626;
array[13071]=30'd900139626;
array[13072]=30'd900139626;
array[13073]=30'd900139626;
array[13074]=30'd900139626;
array[13075]=30'd900139626;
array[13076]=30'd900139626;
array[13077]=30'd900139626;
array[13078]=30'd900139626;
array[13079]=30'd900139626;
array[13080]=30'd900139626;
array[13081]=30'd900139626;
array[13082]=30'd900139626;
array[13083]=30'd873911932;
array[13084]=30'd900139626;
array[13085]=30'd900139626;
array[13086]=30'd900139626;
array[13087]=30'd900139626;
array[13088]=30'd900139626;
array[13089]=30'd900139626;
array[13090]=30'd900139626;
array[13091]=30'd900139626;
array[13092]=30'd900139626;
array[13093]=30'd900139626;
array[13094]=30'd873911932;
array[13095]=30'd873911932;
array[13096]=30'd873911932;
array[13097]=30'd873911932;
array[13098]=30'd527847013;
array[13099]=30'd427157133;
array[13100]=30'd644165300;
array[13101]=30'd653646508;
array[13102]=30'd474371718;
array[13103]=30'd740728401;
array[13104]=30'd941029952;
array[13105]=30'd959928886;
array[13106]=30'd959928886;
array[13107]=30'd959928886;
array[13108]=30'd959928886;
array[13109]=30'd959928886;
array[13110]=30'd959928886;
array[13111]=30'd959928886;
array[13112]=30'd959928886;
array[13113]=30'd959928886;
array[13114]=30'd985089582;
array[13115]=30'd959928886;
array[13116]=30'd959928886;
array[13117]=30'd959928886;
array[13118]=30'd959928886;
array[13119]=30'd959928886;
array[13120]=30'd959928886;
array[13121]=30'd959928886;
array[13122]=30'd959928886;
array[13123]=30'd959928886;
array[13124]=30'd959928886;
array[13125]=30'd941029952;
array[13126]=30'd625391195;
array[13127]=30'd581297788;
array[13128]=30'd549823127;
array[13129]=30'd557159098;
array[13130]=30'd596983478;
array[13131]=30'd452327079;
array[13132]=30'd397801110;
array[13133]=30'd609598119;
array[13134]=30'd609598119;
array[13135]=30'd684081775;
array[13136]=30'd887567935;
array[13137]=30'd778567150;
array[13138]=30'd832058842;
array[13139]=30'd1019742694;
array[13140]=30'd950544914;
array[13141]=30'd785935846;
array[13142]=30'd764964292;
array[13143]=30'd945318330;
array[13144]=30'd1000883648;
array[13145]=30'd945318330;
array[13146]=30'd869807552;
array[13147]=30'd782796193;
array[13148]=30'd888658404;
array[13149]=30'd890710541;
array[13150]=30'd867617357;
array[13151]=30'd873911932;
array[13152]=30'd875034136;
array[13153]=30'd855119352;
array[13154]=30'd855119352;
array[13155]=30'd890710541;
array[13156]=30'd916923947;
array[13157]=30'd900139626;
array[13158]=30'd900139626;
array[13159]=30'd900139626;
array[13160]=30'd900139626;
array[13161]=30'd900139626;
array[13162]=30'd900139626;
array[13163]=30'd900139626;
array[13164]=30'd900139626;
array[13165]=30'd900139626;
array[13166]=30'd900139626;
array[13167]=30'd900139626;
array[13168]=30'd900139626;
array[13169]=30'd900139626;
array[13170]=30'd900139626;
array[13171]=30'd900139626;
array[13172]=30'd900139626;
array[13173]=30'd900139626;
array[13174]=30'd900139626;
array[13175]=30'd900139626;
array[13176]=30'd900139626;
array[13177]=30'd900139626;
array[13178]=30'd900139626;
array[13179]=30'd900139626;
array[13180]=30'd900139626;
array[13181]=30'd900139626;
array[13182]=30'd900139626;
array[13183]=30'd900139626;
array[13184]=30'd900139626;
array[13185]=30'd887567935;
array[13186]=30'd887567935;
array[13187]=30'd887567935;
array[13188]=30'd887567935;
array[13189]=30'd900139626;
array[13190]=30'd900139626;
array[13191]=30'd900139626;
array[13192]=30'd873911932;
array[13193]=30'd873911932;
array[13194]=30'd625391195;
array[13195]=30'd446038641;
array[13196]=30'd644165300;
array[13197]=30'd596983478;
array[13198]=30'd452327079;
array[13199]=30'd433483392;
array[13200]=30'd625391195;
array[13201]=30'd887567935;
array[13202]=30'd959928886;
array[13203]=30'd959928886;
array[13204]=30'd959928886;
array[13205]=30'd959928886;
array[13206]=30'd959928886;
array[13207]=30'd959928886;
array[13208]=30'd959928886;
array[13209]=30'd959928886;
array[13210]=30'd959928886;
array[13211]=30'd959928886;
array[13212]=30'd959928886;
array[13213]=30'd959928886;
array[13214]=30'd959928886;
array[13215]=30'd959928886;
array[13216]=30'd959928886;
array[13217]=30'd959928886;
array[13218]=30'd959928886;
array[13219]=30'd941029952;
array[13220]=30'd887567935;
array[13221]=30'd625391195;
array[13222]=30'd374751849;
array[13223]=30'd636841618;
array[13224]=30'd452327079;
array[13225]=30'd644165300;
array[13226]=30'd549823127;
array[13227]=30'd364251806;
array[13228]=30'd461756049;
array[13229]=30'd636841618;
array[13230]=30'd557159098;
array[13231]=30'd792127082;
array[13232]=30'd887567935;
array[13233]=30'd820526616;
array[13234]=30'd785935846;
array[13235]=30'd904416730;
array[13236]=30'd987238908;
array[13237]=30'd926429685;
array[13238]=30'd764964292;
array[13239]=30'd782796193;
array[13240]=30'd869807552;
array[13241]=30'd906527146;
array[13242]=30'd811098555;
array[13243]=30'd764964292;
array[13244]=30'd870795757;
array[13245]=30'd867617357;
array[13246]=30'd873911932;
array[13247]=30'd873911932;
array[13248]=30'd887567935;
array[13249]=30'd890710541;
array[13250]=30'd910663171;
array[13251]=30'd887567935;
array[13252]=30'd887567935;
array[13253]=30'd900139626;
array[13254]=30'd900139626;
array[13255]=30'd900139626;
array[13256]=30'd873911932;
array[13257]=30'd900139626;
array[13258]=30'd900139626;
array[13259]=30'd900139626;
array[13260]=30'd900139626;
array[13261]=30'd900139626;
array[13262]=30'd900139626;
array[13263]=30'd900139626;
array[13264]=30'd900139626;
array[13265]=30'd900139626;
array[13266]=30'd900139626;
array[13267]=30'd900139626;
array[13268]=30'd900139626;
array[13269]=30'd900139626;
array[13270]=30'd900139626;
array[13271]=30'd900139626;
array[13272]=30'd900139626;
array[13273]=30'd900139626;
array[13274]=30'd900139626;
array[13275]=30'd900139626;
array[13276]=30'd900139626;
array[13277]=30'd900139626;
array[13278]=30'd900139626;
array[13279]=30'd900139626;
array[13280]=30'd887567935;
array[13281]=30'd809995819;
array[13282]=30'd967280137;
array[13283]=30'd875034136;
array[13284]=30'd809995819;
array[13285]=30'd935829023;
array[13286]=30'd887567935;
array[13287]=30'd887567935;
array[13288]=30'd900139626;
array[13289]=30'd900139626;
array[13290]=30'd709314133;
array[13291]=30'd486913656;
array[13292]=30'd636841618;
array[13293]=30'd557159098;
array[13294]=30'd452327079;
array[13295]=30'd427157133;
array[13296]=30'd374751849;
array[13297]=30'd453416554;
array[13298]=30'd709314133;
array[13299]=30'd916923947;
array[13300]=30'd959928886;
array[13301]=30'd959928886;
array[13302]=30'd959928886;
array[13303]=30'd959928886;
array[13304]=30'd959928886;
array[13305]=30'd959928886;
array[13306]=30'd959928886;
array[13307]=30'd959928886;
array[13308]=30'd959928886;
array[13309]=30'd959928886;
array[13310]=30'd959928886;
array[13311]=30'd959928886;
array[13312]=30'd959928886;
array[13313]=30'd959928886;
array[13314]=30'd941029952;
array[13315]=30'd757545539;
array[13316]=30'd455516734;
array[13317]=30'd404111966;
array[13318]=30'd446038641;
array[13319]=30'd581297788;
array[13320]=30'd515208870;
array[13321]=30'd596983478;
array[13322]=30'd427157133;
array[13323]=30'd328601227;
array[13324]=30'd503733877;
array[13325]=30'd636841618;
array[13326]=30'd549823127;
array[13327]=30'd852917899;
array[13328]=30'd900139626;
array[13329]=30'd857219651;
array[13330]=30'd820526616;
array[13331]=30'd832058842;
array[13332]=30'd964180446;
array[13333]=30'd987238908;
array[13334]=30'd855119352;
array[13335]=30'd785935846;
array[13336]=30'd764964292;
array[13337]=30'd764964292;
array[13338]=30'd794289609;
array[13339]=30'd832058842;
array[13340]=30'd890710541;
array[13341]=30'd867617357;
array[13342]=30'd900139626;
array[13343]=30'd873911932;
array[13344]=30'd900139626;
array[13345]=30'd900139626;
array[13346]=30'd900139626;
array[13347]=30'd900139626;
array[13348]=30'd900139626;
array[13349]=30'd900139626;
array[13350]=30'd900139626;
array[13351]=30'd900139626;
array[13352]=30'd900139626;
array[13353]=30'd873911932;
array[13354]=30'd900139626;
array[13355]=30'd900139626;
array[13356]=30'd900139626;
array[13357]=30'd900139626;
array[13358]=30'd900139626;
array[13359]=30'd900139626;
array[13360]=30'd900139626;
array[13361]=30'd900139626;
array[13362]=30'd900139626;
array[13363]=30'd900139626;
array[13364]=30'd900139626;
array[13365]=30'd900139626;
array[13366]=30'd900139626;
array[13367]=30'd900139626;
array[13368]=30'd900139626;
array[13369]=30'd900139626;
array[13370]=30'd900139626;
array[13371]=30'd900139626;
array[13372]=30'd900139626;
array[13373]=30'd900139626;
array[13374]=30'd900139626;
array[13375]=30'd921150041;
array[13376]=30'd898098744;
array[13377]=30'd820526616;
array[13378]=30'd967280137;
array[13379]=30'd855119352;
array[13380]=30'd855119352;
array[13381]=30'd967280137;
array[13382]=30'd875034136;
array[13383]=30'd809995819;
array[13384]=30'd862402083;
array[13385]=30'd887567935;
array[13386]=30'd740728401;
array[13387]=30'd503733877;
array[13388]=30'd636841618;
array[13389]=30'd557159098;
array[13390]=30'd452327079;
array[13391]=30'd427157133;
array[13392]=30'd351684214;
array[13393]=30'd453416554;
array[13394]=30'd404111966;
array[13395]=30'd417793613;
array[13396]=30'd625391195;
array[13397]=30'd794232376;
array[13398]=30'd916923947;
array[13399]=30'd941029952;
array[13400]=30'd959928886;
array[13401]=30'd959928886;
array[13402]=30'd959928886;
array[13403]=30'd959928886;
array[13404]=30'd959928886;
array[13405]=30'd985089582;
array[13406]=30'd959928886;
array[13407]=30'd959928886;
array[13408]=30'd887567935;
array[13409]=30'd794232376;
array[13410]=30'd511088198;
array[13411]=30'd417793613;
array[13412]=30'd453416554;
array[13413]=30'd404111966;
array[13414]=30'd503733877;
array[13415]=30'd461756049;
array[13416]=30'd609598119;
array[13417]=30'd522581659;
array[13418]=30'd300284569;
array[13419]=30'd266734242;
array[13420]=30'd486913656;
array[13421]=30'd636841618;
array[13422]=30'd560346760;
array[13423]=30'd873911932;
array[13424]=30'd900139626;
array[13425]=30'd887567935;
array[13426]=30'd875034136;
array[13427]=30'd785935846;
array[13428]=30'd832058842;
array[13429]=30'd987238908;
array[13430]=30'd950544914;
array[13431]=30'd875034136;
array[13432]=30'd875034136;
array[13433]=30'd855119352;
array[13434]=30'd910663171;
array[13435]=30'd916923947;
array[13436]=30'd887567935;
array[13437]=30'd900139626;
array[13438]=30'd873911932;
array[13439]=30'd873911932;
array[13440]=30'd900139626;
array[13441]=30'd900139626;
array[13442]=30'd900139626;
array[13443]=30'd900139626;
array[13444]=30'd900139626;
array[13445]=30'd900139626;
array[13446]=30'd900139626;
array[13447]=30'd900139626;
array[13448]=30'd900139626;
array[13449]=30'd900139626;
array[13450]=30'd900139626;
array[13451]=30'd900139626;
array[13452]=30'd900139626;
array[13453]=30'd900139626;
array[13454]=30'd900139626;
array[13455]=30'd900139626;
array[13456]=30'd900139626;
array[13457]=30'd900139626;
array[13458]=30'd900139626;
array[13459]=30'd900139626;
array[13460]=30'd900139626;
array[13461]=30'd900139626;
array[13462]=30'd900139626;
array[13463]=30'd900139626;
array[13464]=30'd900139626;
array[13465]=30'd900139626;
array[13466]=30'd900139626;
array[13467]=30'd900139626;
array[13468]=30'd900139626;
array[13469]=30'd900139626;
array[13470]=30'd900139626;
array[13471]=30'd900139626;
array[13472]=30'd921150041;
array[13473]=30'd898098744;
array[13474]=30'd967280137;
array[13475]=30'd875034136;
array[13476]=30'd926429685;
array[13477]=30'd967280137;
array[13478]=30'd844591615;
array[13479]=30'd910663171;
array[13480]=30'd935829023;
array[13481]=30'd887567935;
array[13482]=30'd740735615;
array[13483]=30'd560346760;
array[13484]=30'd636841618;
array[13485]=30'd549823127;
array[13486]=30'd452327079;
array[13487]=30'd433483392;
array[13488]=30'd404111966;
array[13489]=30'd433483392;
array[13490]=30'd410428039;
array[13491]=30'd404111966;
array[13492]=30'd453416554;
array[13493]=30'd404111966;
array[13494]=30'd417793613;
array[13495]=30'd511088198;
array[13496]=30'd666281541;
array[13497]=30'd794232376;
array[13498]=30'd840392271;
array[13499]=30'd867617357;
array[13500]=30'd867617357;
array[13501]=30'd794232376;
array[13502]=30'd709314133;
array[13503]=30'd666281541;
array[13504]=30'd679964212;
array[13505]=30'd757545539;
array[13506]=30'd334932558;
array[13507]=30'd455516734;
array[13508]=30'd453416554;
array[13509]=30'd364251806;
array[13510]=30'd522581659;
array[13511]=30'd522581659;
array[13512]=30'd549823127;
array[13513]=30'd364251806;
array[13514]=30'd266734242;
array[13515]=30'd351684214;
array[13516]=30'd522581659;
array[13517]=30'd636841618;
array[13518]=30'd581297788;
array[13519]=30'd873911932;
array[13520]=30'd900139626;
array[13521]=30'd900139626;
array[13522]=30'd898098744;
array[13523]=30'd857219651;
array[13524]=30'd785935846;
array[13525]=30'd888658404;
array[13526]=30'd1019742694;
array[13527]=30'd987238908;
array[13528]=30'd950544914;
array[13529]=30'd950544914;
array[13530]=30'd967280137;
array[13531]=30'd941029952;
array[13532]=30'd900139626;
array[13533]=30'd900139626;
array[13534]=30'd873911932;
array[13535]=30'd900139626;
array[13536]=30'd900139626;
array[13537]=30'd900139626;
array[13538]=30'd900139626;
array[13539]=30'd900139626;
array[13540]=30'd900139626;
array[13541]=30'd900139626;
array[13542]=30'd921150041;
array[13543]=30'd898098744;
array[13544]=30'd875034136;
array[13545]=30'd844591615;
array[13546]=30'd820526616;
array[13547]=30'd898098744;
array[13548]=30'd887567935;
array[13549]=30'd887567935;
array[13550]=30'd900139626;
array[13551]=30'd900139626;
array[13552]=30'd900139626;
array[13553]=30'd900139626;
array[13554]=30'd900139626;
array[13555]=30'd900139626;
array[13556]=30'd900139626;
array[13557]=30'd900139626;
array[13558]=30'd900139626;
array[13559]=30'd900139626;
array[13560]=30'd900139626;
array[13561]=30'd900139626;
array[13562]=30'd900139626;
array[13563]=30'd900139626;
array[13564]=30'd900139626;
array[13565]=30'd900139626;
array[13566]=30'd900139626;
array[13567]=30'd900139626;
array[13568]=30'd921150041;
array[13569]=30'd898098744;
array[13570]=30'd875034136;
array[13571]=30'd875034136;
array[13572]=30'd910663171;
array[13573]=30'd888658404;
array[13574]=30'd855119352;
array[13575]=30'd967280137;
array[13576]=30'd916923947;
array[13577]=30'd867617357;
array[13578]=30'd740735615;
array[13579]=30'd581297788;
array[13580]=30'd644165300;
array[13581]=30'd485848753;
array[13582]=30'd461756049;
array[13583]=30'd404111966;
array[13584]=30'd410428039;
array[13585]=30'd433483392;
array[13586]=30'd364251806;
array[13587]=30'd351684214;
array[13588]=30'd446038641;
array[13589]=30'd446038641;
array[13590]=30'd433483392;
array[13591]=30'd453416554;
array[13592]=30'd404111966;
array[13593]=30'd455516734;
array[13594]=30'd794232376;
array[13595]=30'd794232376;
array[13596]=30'd794232376;
array[13597]=30'd794232376;
array[13598]=30'd792127082;
array[13599]=30'd792127082;
array[13600]=30'd821480030;
array[13601]=30'd757545539;
array[13602]=30'd245885528;
array[13603]=30'd312961612;
array[13604]=30'd404111966;
array[13605]=30'd446038641;
array[13606]=30'd461756049;
array[13607]=30'd557159098;
array[13608]=30'd452327079;
array[13609]=30'd266734242;
array[13610]=30'd364251806;
array[13611]=30'd351684214;
array[13612]=30'd522581659;
array[13613]=30'd609598119;
array[13614]=30'd625391195;
array[13615]=30'd900139626;
array[13616]=30'd900139626;
array[13617]=30'd873911932;
array[13618]=30'd900139626;
array[13619]=30'd898098744;
array[13620]=30'd820526616;
array[13621]=30'd778567150;
array[13622]=30'd869807552;
array[13623]=30'd849905057;
array[13624]=30'd811098555;
array[13625]=30'd811098555;
array[13626]=30'd888658404;
array[13627]=30'd916923947;
array[13628]=30'd900139626;
array[13629]=30'd873911932;
array[13630]=30'd873911932;
array[13631]=30'd873911932;
array[13632]=30'd900139626;
array[13633]=30'd900139626;
array[13634]=30'd900139626;
array[13635]=30'd900139626;
array[13636]=30'd900139626;
array[13637]=30'd900139626;
array[13638]=30'd875034136;
array[13639]=30'd785935846;
array[13640]=30'd832058842;
array[13641]=30'd869807552;
array[13642]=30'd832058842;
array[13643]=30'd778567150;
array[13644]=30'd844591615;
array[13645]=30'd890710541;
array[13646]=30'd887567935;
array[13647]=30'd900139626;
array[13648]=30'd921150041;
array[13649]=30'd921150041;
array[13650]=30'd898098744;
array[13651]=30'd887567935;
array[13652]=30'd887567935;
array[13653]=30'd900139626;
array[13654]=30'd900139626;
array[13655]=30'd900139626;
array[13656]=30'd900139626;
array[13657]=30'd900139626;
array[13658]=30'd900139626;
array[13659]=30'd900139626;
array[13660]=30'd900139626;
array[13661]=30'd900139626;
array[13662]=30'd921150041;
array[13663]=30'd898098744;
array[13664]=30'd875034136;
array[13665]=30'd820526616;
array[13666]=30'd855119352;
array[13667]=30'd832058842;
array[13668]=30'd785935846;
array[13669]=30'd820487650;
array[13670]=30'd888658404;
array[13671]=30'd910663171;
array[13672]=30'd887567935;
array[13673]=30'd900139626;
array[13674]=30'd709304966;
array[13675]=30'd636841618;
array[13676]=30'd644165300;
array[13677]=30'd485848753;
array[13678]=30'd427157133;
array[13679]=30'd334965361;
array[13680]=30'd404111966;
array[13681]=30'd446038641;
array[13682]=30'd410428039;
array[13683]=30'd278304367;
array[13684]=30'd446038641;
array[13685]=30'd427157133;
array[13686]=30'd427157133;
array[13687]=30'd433483392;
array[13688]=30'd334965361;
array[13689]=30'd352820791;
array[13690]=30'd821480030;
array[13691]=30'd821480030;
array[13692]=30'd821480030;
array[13693]=30'd821480030;
array[13694]=30'd821480030;
array[13695]=30'd821480030;
array[13696]=30'd679964212;
array[13697]=30'd393770575;
array[13698]=30'd274187850;
array[13699]=30'd274187850;
array[13700]=30'd259444308;
array[13701]=30'd446038641;
array[13702]=30'd549823127;
array[13703]=30'd515208870;
array[13704]=30'd364251806;
array[13705]=30'd334965361;
array[13706]=30'd404111966;
array[13707]=30'd374751849;
array[13708]=30'd522581659;
array[13709]=30'd609598119;
array[13710]=30'd684081775;
array[13711]=30'd900139626;
array[13712]=30'd900139626;
array[13713]=30'd873911932;
array[13714]=30'd900139626;
array[13715]=30'd900139626;
array[13716]=30'd898098744;
array[13717]=30'd820526616;
array[13718]=30'd785935846;
array[13719]=30'd794289609;
array[13720]=30'd794289609;
array[13721]=30'd820487650;
array[13722]=30'd844591615;
array[13723]=30'd887567935;
array[13724]=30'd900139626;
array[13725]=30'd900139626;
array[13726]=30'd873911932;
array[13727]=30'd873911932;
array[13728]=30'd900139626;
array[13729]=30'd900139626;
array[13730]=30'd900139626;
array[13731]=30'd900139626;
array[13732]=30'd900139626;
array[13733]=30'd921150041;
array[13734]=30'd875034136;
array[13735]=30'd904416730;
array[13736]=30'd964180446;
array[13737]=30'd987238908;
array[13738]=30'd987238908;
array[13739]=30'd926429685;
array[13740]=30'd794289609;
array[13741]=30'd820487650;
array[13742]=30'd890710541;
array[13743]=30'd887567935;
array[13744]=30'd898098744;
array[13745]=30'd820526616;
array[13746]=30'd778567150;
array[13747]=30'd844591615;
array[13748]=30'd887567935;
array[13749]=30'd900139626;
array[13750]=30'd900139626;
array[13751]=30'd900139626;
array[13752]=30'd900139626;
array[13753]=30'd900139626;
array[13754]=30'd900139626;
array[13755]=30'd900139626;
array[13756]=30'd900139626;
array[13757]=30'd921150041;
array[13758]=30'd921150041;
array[13759]=30'd820526616;
array[13760]=30'd875034136;
array[13761]=30'd987238908;
array[13762]=30'd964180446;
array[13763]=30'd926429685;
array[13764]=30'd926429685;
array[13765]=30'd888658404;
array[13766]=30'd820487650;
array[13767]=30'd935829023;
array[13768]=30'd887567935;
array[13769]=30'd900139626;
array[13770]=30'd684081775;
array[13771]=30'd626373227;
array[13772]=30'd609598119;
array[13773]=30'd452327079;
array[13774]=30'd328601227;
array[13775]=30'd305565277;
array[13776]=30'd374751849;
array[13777]=30'd446038641;
array[13778]=30'd410428039;
array[13779]=30'd259444308;
array[13780]=30'd446038641;
array[13781]=30'd446038641;
array[13782]=30'd433483392;
array[13783]=30'd404111966;
array[13784]=30'd274187850;
array[13785]=30'd352820791;
array[13786]=30'd757545539;
array[13787]=30'd821480030;
array[13788]=30'd821480030;
array[13789]=30'd792127082;
array[13790]=30'd709314133;
array[13791]=30'd472349226;
array[13792]=30'd274187850;
array[13793]=30'd302559805;
array[13794]=30'd302559805;
array[13795]=30'd302559805;
array[13796]=30'd334932558;
array[13797]=30'd446038641;
array[13798]=30'd549823127;
array[13799]=30'd427157133;
array[13800]=30'd266734242;
array[13801]=30'd404111966;
array[13802]=30'd351684214;
array[13803]=30'd374751849;
array[13804]=30'd496374434;
array[13805]=30'd549823127;
array[13806]=30'd709304966;
array[13807]=30'd900139626;
array[13808]=30'd873911932;
array[13809]=30'd873911932;
array[13810]=30'd900139626;
array[13811]=30'd873911932;
array[13812]=30'd900139626;
array[13813]=30'd887567935;
array[13814]=30'd887567935;
array[13815]=30'd887567935;
array[13816]=30'd887567935;
array[13817]=30'd887567935;
array[13818]=30'd887567935;
array[13819]=30'd900139626;
array[13820]=30'd900139626;
array[13821]=30'd873911932;
array[13822]=30'd873911932;
array[13823]=30'd873911932;
array[13824]=30'd900139626;
array[13825]=30'd900139626;
array[13826]=30'd900139626;
array[13827]=30'd900139626;
array[13828]=30'd900139626;
array[13829]=30'd921150041;
array[13830]=30'd967280137;
array[13831]=30'd742923790;
array[13832]=30'd778567150;
array[13833]=30'd875034136;
array[13834]=30'd950544914;
array[13835]=30'd987238908;
array[13836]=30'd964180446;
array[13837]=30'd832058842;
array[13838]=30'd820487650;
array[13839]=30'd890710541;
array[13840]=30'd898098744;
array[13841]=30'd875034136;
array[13842]=30'd946320871;
array[13843]=30'd910663171;
array[13844]=30'd887567935;
array[13845]=30'd900139626;
array[13846]=30'd900139626;
array[13847]=30'd900139626;
array[13848]=30'd900139626;
array[13849]=30'd900139626;
array[13850]=30'd900139626;
array[13851]=30'd900139626;
array[13852]=30'd900139626;
array[13853]=30'd921150041;
array[13854]=30'd857219651;
array[13855]=30'd855119352;
array[13856]=30'd1019742694;
array[13857]=30'd926429685;
array[13858]=30'd855119352;
array[13859]=30'd832058842;
array[13860]=30'd832058842;
array[13861]=30'd869807552;
array[13862]=30'd832058842;
array[13863]=30'd910663171;
array[13864]=30'd916923947;
array[13865]=30'd900139626;
array[13866]=30'd625391195;
array[13867]=30'd636841618;
array[13868]=30'd609598119;
array[13869]=30'd427157133;
array[13870]=30'd351684214;
array[13871]=30'd334965361;
array[13872]=30'd351684214;
array[13873]=30'd446038641;
array[13874]=30'd453416554;
array[13875]=30'd259444308;
array[13876]=30'd446038641;
array[13877]=30'd446038641;
array[13878]=30'd384241245;
array[13879]=30'd294104668;
array[13880]=30'd302559805;
array[13881]=30'd393770575;
array[13882]=30'd709314133;
array[13883]=30'd821480030;
array[13884]=30'd792127082;
array[13885]=30'd593947240;
array[13886]=30'd294104668;
array[13887]=30'd302559805;
array[13888]=30'd281613891;
array[13889]=30'd281613891;
array[13890]=30'd302559805;
array[13891]=30'd302559805;
array[13892]=30'd334932558;
array[13893]=30'd560346760;
array[13894]=30'd461756049;
array[13895]=30'd364251806;
array[13896]=30'd278304367;
array[13897]=30'd410428039;
array[13898]=30'd305565277;
array[13899]=30'd404111966;
array[13900]=30'd461756049;
array[13901]=30'd549823127;
array[13902]=30'd740735615;
array[13903]=30'd900139626;
array[13904]=30'd873911932;
array[13905]=30'd873911932;
array[13906]=30'd873911932;
array[13907]=30'd873911932;
array[13908]=30'd900139626;
array[13909]=30'd900139626;
array[13910]=30'd900139626;
array[13911]=30'd900139626;
array[13912]=30'd900139626;
array[13913]=30'd900139626;
array[13914]=30'd900139626;
array[13915]=30'd900139626;
array[13916]=30'd900139626;
array[13917]=30'd873911932;
array[13918]=30'd873911932;
array[13919]=30'd873911932;
array[13920]=30'd900139626;
array[13921]=30'd900139626;
array[13922]=30'd900139626;
array[13923]=30'd900139626;
array[13924]=30'd900139626;
array[13925]=30'd840392271;
array[13926]=30'd742923790;
array[13927]=30'd519570948;
array[13928]=30'd708323812;
array[13929]=30'd785935846;
array[13930]=30'd785935846;
array[13931]=30'd888658404;
array[13932]=30'd964180446;
array[13933]=30'd964180446;
array[13934]=30'd794289609;
array[13935]=30'd888658404;
array[13936]=30'd935829023;
array[13937]=30'd950544914;
array[13938]=30'd967280137;
array[13939]=30'd916923947;
array[13940]=30'd887567935;
array[13941]=30'd900139626;
array[13942]=30'd900139626;
array[13943]=30'd900139626;
array[13944]=30'd900139626;
array[13945]=30'd900139626;
array[13946]=30'd900139626;
array[13947]=30'd900139626;
array[13948]=30'd921150041;
array[13949]=30'd857219651;
array[13950]=30'd855119352;
array[13951]=30'd964180446;
array[13952]=30'd904416730;
array[13953]=30'd785935846;
array[13954]=30'd832058842;
array[13955]=30'd904416730;
array[13956]=30'd869807552;
array[13957]=30'd869807552;
array[13958]=30'd869807552;
array[13959]=30'd888658404;
array[13960]=30'd916923947;
array[13961]=30'd900139626;
array[13962]=30'd593947240;
array[13963]=30'd636841618;
array[13964]=30'd557159098;
array[13965]=30'd397801110;
array[13966]=30'd351684214;
array[13967]=30'd374751849;
array[13968]=30'd334932558;
array[13969]=30'd446038641;
array[13970]=30'd453416554;
array[13971]=30'd334932558;
array[13972]=30'd361192034;
array[13973]=30'd312961612;
array[13974]=30'd274187850;
array[13975]=30'd302559805;
array[13976]=30'd302559805;
array[13977]=30'd393770575;
array[13978]=30'd778555959;
array[13979]=30'd778555959;
array[13980]=30'd506984008;
array[13981]=30'd274187850;
array[13982]=30'd302559805;
array[13983]=30'd281613891;
array[13984]=30'd281613891;
array[13985]=30'd281613891;
array[13986]=30'd281613891;
array[13987]=30'd274187850;
array[13988]=30'd453416554;
array[13989]=30'd522581659;
array[13990]=30'd427157133;
array[13991]=30'd278304367;
array[13992]=30'd384241245;
array[13993]=30'd417793613;
array[13994]=30'd305565277;
array[13995]=30'd404111966;
array[13996]=30'd461756049;
array[13997]=30'd522581659;
array[13998]=30'd792127082;
array[13999]=30'd900139626;
array[14000]=30'd873911932;
array[14001]=30'd873911932;
array[14002]=30'd900139626;
array[14003]=30'd900139626;
array[14004]=30'd900139626;
array[14005]=30'd873911932;
array[14006]=30'd873911932;
array[14007]=30'd900139626;
array[14008]=30'd900139626;
array[14009]=30'd900139626;
array[14010]=30'd900139626;
array[14011]=30'd873911932;
array[14012]=30'd873911932;
array[14013]=30'd900139626;
array[14014]=30'd900139626;
array[14015]=30'd900139626;
array[14016]=30'd900139626;
array[14017]=30'd900139626;
array[14018]=30'd900139626;
array[14019]=30'd900139626;
array[14020]=30'd804758111;
array[14021]=30'd655912516;
array[14022]=30'd651672075;
array[14023]=30'd778567150;
array[14024]=30'd752351692;
array[14025]=30'd904416730;
array[14026]=30'd869807552;
array[14027]=30'd811098555;
array[14028]=30'd910663171;
array[14029]=30'd987238908;
array[14030]=30'd832058842;
array[14031]=30'd832058842;
array[14032]=30'd910663171;
array[14033]=30'd855119352;
array[14034]=30'd820487650;
array[14035]=30'd844591615;
array[14036]=30'd890710541;
array[14037]=30'd900139626;
array[14038]=30'd900139626;
array[14039]=30'd900139626;
array[14040]=30'd900139626;
array[14041]=30'd900139626;
array[14042]=30'd900139626;
array[14043]=30'd900139626;
array[14044]=30'd921150041;
array[14045]=30'd875034136;
array[14046]=30'd964180446;
array[14047]=30'd964180446;
array[14048]=30'd785935846;
array[14049]=30'd904416730;
array[14050]=30'd904416730;
array[14051]=30'd945318330;
array[14052]=30'd849905057;
array[14053]=30'd811098555;
array[14054]=30'd906527146;
array[14055]=30'd869807552;
array[14056]=30'd916923947;
array[14057]=30'd900139626;
array[14058]=30'd571937394;
array[14059]=30'd636841618;
array[14060]=30'd549823127;
array[14061]=30'd364251806;
array[14062]=30'd305565277;
array[14063]=30'd404111966;
array[14064]=30'd361192034;
array[14065]=30'd334965361;
array[14066]=30'd361192034;
array[14067]=30'd245885528;
array[14068]=30'd245885528;
array[14069]=30'd238603832;
array[14070]=30'd253299274;
array[14071]=30'd302559805;
array[14072]=30'd281613891;
array[14073]=30'd302559805;
array[14074]=30'd733487691;
array[14075]=30'd431516230;
array[14076]=30'd238603832;
array[14077]=30'd302559805;
array[14078]=30'd281613891;
array[14079]=30'd281613891;
array[14080]=30'd281613891;
array[14081]=30'd281613891;
array[14082]=30'd253299274;
array[14083]=30'd274187850;
array[14084]=30'd560346760;
array[14085]=30'd461756049;
array[14086]=30'd364251806;
array[14087]=30'd232189540;
array[14088]=30'd305565277;
array[14089]=30'd361192034;
array[14090]=30'd305565277;
array[14091]=30'd374751849;
array[14092]=30'd486913656;
array[14093]=30'd522581659;
array[14094]=30'd821480030;
array[14095]=30'd900139626;
array[14096]=30'd900139626;
array[14097]=30'd900139626;
array[14098]=30'd900139626;
array[14099]=30'd900139626;
array[14100]=30'd900139626;
array[14101]=30'd873911932;
array[14102]=30'd900139626;
array[14103]=30'd900139626;
array[14104]=30'd900139626;
array[14105]=30'd900139626;
array[14106]=30'd900139626;
array[14107]=30'd900139626;
array[14108]=30'd900139626;
array[14109]=30'd900139626;
array[14110]=30'd900139626;
array[14111]=30'd900139626;
array[14112]=30'd900139626;
array[14113]=30'd900139626;
array[14114]=30'd900139626;
array[14115]=30'd873911932;
array[14116]=30'd709314133;
array[14117]=30'd820526616;
array[14118]=30'd1033359876;
array[14119]=30'd1033359876;
array[14120]=30'd987238908;
array[14121]=30'd785935846;
array[14122]=30'd869807552;
array[14123]=30'd811098555;
array[14124]=30'd888658404;
array[14125]=30'd926429685;
array[14126]=30'd832058842;
array[14127]=30'd820487650;
array[14128]=30'd910663171;
array[14129]=30'd832058842;
array[14130]=30'd832058842;
array[14131]=30'd820487650;
array[14132]=30'd890710541;
array[14133]=30'd887567935;
array[14134]=30'd900139626;
array[14135]=30'd900139626;
array[14136]=30'd900139626;
array[14137]=30'd900139626;
array[14138]=30'd900139626;
array[14139]=30'd900139626;
array[14140]=30'd921150041;
array[14141]=30'd820526616;
array[14142]=30'd926429685;
array[14143]=30'd926429685;
array[14144]=30'd832058842;
array[14145]=30'd945318330;
array[14146]=30'd811098555;
array[14147]=30'd811098555;
array[14148]=30'd833137031;
array[14149]=30'd833137031;
array[14150]=30'd811098555;
array[14151]=30'd929554891;
array[14152]=30'd916923947;
array[14153]=30'd900139626;
array[14154]=30'd527847013;
array[14155]=30'd636841618;
array[14156]=30'd549823127;
array[14157]=30'd351684214;
array[14158]=30'd278304367;
array[14159]=30'd361192034;
array[14160]=30'd393770575;
array[14161]=30'd451435107;
array[14162]=30'd453527098;
array[14163]=30'd361277993;
array[14164]=30'd281613891;
array[14165]=30'd238603832;
array[14166]=30'd281613891;
array[14167]=30'd281613891;
array[14168]=30'd281613891;
array[14169]=30'd253299274;
array[14170]=30'd302559805;
array[14171]=30'd253299274;
array[14172]=30'd302559805;
array[14173]=30'd281613891;
array[14174]=30'd281613891;
array[14175]=30'd281613891;
array[14176]=30'd281613891;
array[14177]=30'd281613891;
array[14178]=30'd238603832;
array[14179]=30'd482780758;
array[14180]=30'd503733877;
array[14181]=30'd427157133;
array[14182]=30'd305565277;
array[14183]=30'd232189540;
array[14184]=30'd274187850;
array[14185]=30'd274187850;
array[14186]=30'd219656764;
array[14187]=30'd334932558;
array[14188]=30'd446038641;
array[14189]=30'd503733877;
array[14190]=30'd792127082;
array[14191]=30'd900139626;
array[14192]=30'd873911932;
array[14193]=30'd900139626;
array[14194]=30'd900139626;
array[14195]=30'd900139626;
array[14196]=30'd900139626;
array[14197]=30'd900139626;
array[14198]=30'd900139626;
array[14199]=30'd900139626;
array[14200]=30'd900139626;
array[14201]=30'd900139626;
array[14202]=30'd900139626;
array[14203]=30'd900139626;
array[14204]=30'd900139626;
array[14205]=30'd900139626;
array[14206]=30'd900139626;
array[14207]=30'd900139626;
array[14208]=30'd900139626;
array[14209]=30'd900139626;
array[14210]=30'd900139626;
array[14211]=30'd747092585;
array[14212]=30'd573005379;
array[14213]=30'd935829023;
array[14214]=30'd1033359876;
array[14215]=30'd1033359876;
array[14216]=30'd1033359876;
array[14217]=30'd987238908;
array[14218]=30'd778567150;
array[14219]=30'd869807552;
array[14220]=30'd820487650;
array[14221]=30'd926429685;
array[14222]=30'd855119352;
array[14223]=30'd832058842;
array[14224]=30'd946320871;
array[14225]=30'd987238908;
array[14226]=30'd1019742694;
array[14227]=30'd967280137;
array[14228]=30'd916923947;
array[14229]=30'd887567935;
array[14230]=30'd900139626;
array[14231]=30'd900139626;
array[14232]=30'd900139626;
array[14233]=30'd900139626;
array[14234]=30'd900139626;
array[14235]=30'd900139626;
array[14236]=30'd921150041;
array[14237]=30'd898098744;
array[14238]=30'd875034136;
array[14239]=30'd926429685;
array[14240]=30'd785935846;
array[14241]=30'd869807552;
array[14242]=30'd869807552;
array[14243]=30'd906527146;
array[14244]=30'd849905057;
array[14245]=30'd869807552;
array[14246]=30'd929554891;
array[14247]=30'd910663171;
array[14248]=30'd887567935;
array[14249]=30'd900139626;
array[14250]=30'd527847013;
array[14251]=30'd636841618;
array[14252]=30'd522581659;
array[14253]=30'd278304367;
array[14254]=30'd339237463;
array[14255]=30'd483946067;
array[14256]=30'd487155275;
array[14257]=30'd472478290;
array[14258]=30'd472478290;
array[14259]=30'd412701256;
array[14260]=30'd281613891;
array[14261]=30'd253299274;
array[14262]=30'd281613891;
array[14263]=30'd281613891;
array[14264]=30'd281613891;
array[14265]=30'd253299274;
array[14266]=30'd253299274;
array[14267]=30'd302559805;
array[14268]=30'd281613891;
array[14269]=30'd281613891;
array[14270]=30'd281613891;
array[14271]=30'd281613891;
array[14272]=30'd281613891;
array[14273]=30'd302559805;
array[14274]=30'd312961612;
array[14275]=30'd553016910;
array[14276]=30'd427157133;
array[14277]=30'd364251806;
array[14278]=30'd294104668;
array[14279]=30'd274187850;
array[14280]=30'd339237463;
array[14281]=30'd356077132;
array[14282]=30'd431516230;
array[14283]=30'd393770575;
array[14284]=30'd384241245;
array[14285]=30'd527847013;
array[14286]=30'd740735615;
array[14287]=30'd900139626;
array[14288]=30'd900139626;
array[14289]=30'd900139626;
array[14290]=30'd900139626;
array[14291]=30'd900139626;
array[14292]=30'd900139626;
array[14293]=30'd900139626;
array[14294]=30'd900139626;
array[14295]=30'd900139626;
array[14296]=30'd900139626;
array[14297]=30'd900139626;
array[14298]=30'd900139626;
array[14299]=30'd900139626;
array[14300]=30'd900139626;
array[14301]=30'd900139626;
array[14302]=30'd900139626;
array[14303]=30'd900139626;
array[14304]=30'd900139626;
array[14305]=30'd900139626;
array[14306]=30'd900139626;
array[14307]=30'd900139626;
array[14308]=30'd840392271;
array[14309]=30'd875034136;
array[14310]=30'd1033359876;
array[14311]=30'd1033359876;
array[14312]=30'd1033359876;
array[14313]=30'd1033359876;
array[14314]=30'd964180446;
array[14315]=30'd752351692;
array[14316]=30'd794289609;
array[14317]=30'd926429685;
array[14318]=30'd869807552;
array[14319]=30'd820487650;
array[14320]=30'd910663171;
array[14321]=30'd926429685;
array[14322]=30'd935829023;
array[14323]=30'd935829023;
array[14324]=30'd916923947;
array[14325]=30'd941029952;
array[14326]=30'd900139626;
array[14327]=30'd900139626;
array[14328]=30'd900139626;
array[14329]=30'd900139626;
array[14330]=30'd900139626;
array[14331]=30'd900139626;
array[14332]=30'd921150041;
array[14333]=30'd921150041;
array[14334]=30'd898098744;
array[14335]=30'd935829023;
array[14336]=30'd875034136;
array[14337]=30'd855119352;
array[14338]=30'd855119352;
array[14339]=30'd888658404;
array[14340]=30'd888658404;
array[14341]=30'd967280137;
array[14342]=30'd935829023;
array[14343]=30'd916923947;
array[14344]=30'd900139626;
array[14345]=30'd900139626;
array[14346]=30'd571937394;
array[14347]=30'd636841618;
array[14348]=30'd496374434;
array[14349]=30'd278304367;
array[14350]=30'd431516230;
array[14351]=30'd518580800;
array[14352]=30'd472478290;
array[14353]=30'd487155275;
array[14354]=30'd487155275;
array[14355]=30'd459884097;
array[14356]=30'd317277759;
array[14357]=30'd253299274;
array[14358]=30'd281613891;
array[14359]=30'd281613891;
array[14360]=30'd281613891;
array[14361]=30'd238603832;
array[14362]=30'd206107200;
array[14363]=30'd281613891;
array[14364]=30'd281613891;
array[14365]=30'd281613891;
array[14366]=30'd281613891;
array[14367]=30'd281613891;
array[14368]=30'd281613891;
array[14369]=30'd238603832;
array[14370]=30'd455516734;
array[14371]=30'd503733877;
array[14372]=30'd427157133;
array[14373]=30'd334965361;
array[14374]=30'd334965361;
array[14375]=30'd431516230;
array[14376]=30'd459884097;
array[14377]=30'd459884097;
array[14378]=30'd459884097;
array[14379]=30'd459884097;
array[14380]=30'd431516230;
array[14381]=30'd361192034;
array[14382]=30'd757545539;
array[14383]=30'd900139626;
array[14384]=30'd900139626;
array[14385]=30'd900139626;
array[14386]=30'd900139626;
array[14387]=30'd900139626;
array[14388]=30'd900139626;
array[14389]=30'd900139626;
array[14390]=30'd900139626;
array[14391]=30'd900139626;
array[14392]=30'd900139626;
array[14393]=30'd900139626;
array[14394]=30'd900139626;
array[14395]=30'd900139626;
array[14396]=30'd900139626;
array[14397]=30'd900139626;
array[14398]=30'd900139626;
array[14399]=30'd900139626;
array[14400]=30'd900139626;
array[14401]=30'd900139626;
array[14402]=30'd900139626;
array[14403]=30'd900139626;
array[14404]=30'd900139626;
array[14405]=30'd778555959;
array[14406]=30'd950544914;
array[14407]=30'd1033359876;
array[14408]=30'd1033359876;
array[14409]=30'd1033359876;
array[14410]=30'd1033359876;
array[14411]=30'd964180446;
array[14412]=30'd778567150;
array[14413]=30'd855119352;
array[14414]=30'd785935846;
array[14415]=30'd888658404;
array[14416]=30'd820487650;
array[14417]=30'd742923790;
array[14418]=30'd757556731;
array[14419]=30'd778555959;
array[14420]=30'd794232376;
array[14421]=30'd840392271;
array[14422]=30'd887567935;
array[14423]=30'd900139626;
array[14424]=30'd900139626;
array[14425]=30'd900139626;
array[14426]=30'd900139626;
array[14427]=30'd921150041;
array[14428]=30'd921150041;
array[14429]=30'd921150041;
array[14430]=30'd921150041;
array[14431]=30'd921150041;
array[14432]=30'd921150041;
array[14433]=30'd921150041;
array[14434]=30'd898098744;
array[14435]=30'd935829023;
array[14436]=30'd935829023;
array[14437]=30'd916923947;
array[14438]=30'd921150041;
array[14439]=30'd900139626;
array[14440]=30'd900139626;
array[14441]=30'd900139626;
array[14442]=30'd593947240;
array[14443]=30'd653676161;
array[14444]=30'd474371718;
array[14445]=30'd294104668;
array[14446]=30'd451435107;
array[14447]=30'd472478290;
array[14448]=30'd487155275;
array[14449]=30'd487155275;
array[14450]=30'd487155275;
array[14451]=30'd472478290;
array[14452]=30'd356077132;
array[14453]=30'd281613891;
array[14454]=30'd281613891;
array[14455]=30'd281613891;
array[14456]=30'd238603832;
array[14457]=30'd253299274;
array[14458]=30'd206107200;
array[14459]=30'd238603832;
array[14460]=30'd281613891;
array[14461]=30'd281613891;
array[14462]=30'd281613891;
array[14463]=30'd281613891;
array[14464]=30'd281613891;
array[14465]=30'd274187850;
array[14466]=30'd527847013;
array[14467]=30'd433483392;
array[14468]=30'd374751849;
array[14469]=30'd351684214;
array[14470]=30'd361192034;
array[14471]=30'd483946067;
array[14472]=30'd472478290;
array[14473]=30'd472478290;
array[14474]=30'd472478290;
array[14475]=30'd472478290;
array[14476]=30'd459884097;
array[14477]=30'd431516230;
array[14478]=30'd617068069;
array[14479]=30'd921150041;
array[14480]=30'd900139626;
array[14481]=30'd900139626;
array[14482]=30'd900139626;
array[14483]=30'd900139626;
array[14484]=30'd900139626;
array[14485]=30'd900139626;
array[14486]=30'd900139626;
array[14487]=30'd900139626;
array[14488]=30'd900139626;
array[14489]=30'd900139626;
array[14490]=30'd900139626;
array[14491]=30'd900139626;
array[14492]=30'd900139626;
array[14493]=30'd900139626;
array[14494]=30'd900139626;
array[14495]=30'd900139626;
array[14496]=30'd900139626;
array[14497]=30'd900139626;
array[14498]=30'd921150041;
array[14499]=30'd900139626;
array[14500]=30'd921150041;
array[14501]=30'd921150041;
array[14502]=30'd857219651;
array[14503]=30'd935829023;
array[14504]=30'd1033359876;
array[14505]=30'd1033359876;
array[14506]=30'd1033359876;
array[14507]=30'd1033359876;
array[14508]=30'd987238908;
array[14509]=30'd708323812;
array[14510]=30'd855119352;
array[14511]=30'd926429685;
array[14512]=30'd757556731;
array[14513]=30'd757556731;
array[14514]=30'd890710541;
array[14515]=30'd887567935;
array[14516]=30'd887567935;
array[14517]=30'd809995819;
array[14518]=30'd757545539;
array[14519]=30'd757545539;
array[14520]=30'd840392271;
array[14521]=30'd887567935;
array[14522]=30'd900139626;
array[14523]=30'd900139626;
array[14524]=30'd921150041;
array[14525]=30'd921150041;
array[14526]=30'd921150041;
array[14527]=30'd921150041;
array[14528]=30'd921150041;
array[14529]=30'd921150041;
array[14530]=30'd921150041;
array[14531]=30'd921150041;
array[14532]=30'd900139626;
array[14533]=30'd900139626;
array[14534]=30'd900139626;
array[14535]=30'd900139626;
array[14536]=30'd900139626;
array[14537]=30'd900139626;
array[14538]=30'd549944915;
array[14539]=30'd626373227;
array[14540]=30'd503733877;
array[14541]=30'd294104668;
array[14542]=30'd483946067;
array[14543]=30'd472478290;
array[14544]=30'd472478290;
array[14545]=30'd487155275;
array[14546]=30'd472478290;
array[14547]=30'd472478290;
array[14548]=30'd412701256;
array[14549]=30'd317277759;
array[14550]=30'd253299274;
array[14551]=30'd238603832;
array[14552]=30'd206107200;
array[14553]=30'd176749120;
array[14554]=30'd238603832;
array[14555]=30'd238603832;
array[14556]=30'd281613891;
array[14557]=30'd281613891;
array[14558]=30'd281613891;
array[14559]=30'd317277759;
array[14560]=30'd378082860;
array[14561]=30'd352820791;
array[14562]=30'd560346760;
array[14563]=30'd410428039;
array[14564]=30'd259444308;
array[14565]=30'd417793613;
array[14566]=30'd339237463;
array[14567]=30'd483946067;
array[14568]=30'd472478290;
array[14569]=30'd472478290;
array[14570]=30'd472478290;
array[14571]=30'd472478290;
array[14572]=30'd459884097;
array[14573]=30'd412701256;
array[14574]=30'd431516230;
array[14575]=30'd804758111;
array[14576]=30'd900139626;
array[14577]=30'd900139626;
array[14578]=30'd900139626;
array[14579]=30'd900139626;
array[14580]=30'd900139626;
array[14581]=30'd900139626;
array[14582]=30'd900139626;
array[14583]=30'd900139626;
array[14584]=30'd900139626;
array[14585]=30'd900139626;
array[14586]=30'd900139626;
array[14587]=30'd900139626;
array[14588]=30'd900139626;
array[14589]=30'd900139626;
array[14590]=30'd900139626;
array[14591]=30'd900139626;
array[14592]=30'd900139626;
array[14593]=30'd900139626;
array[14594]=30'd900139626;
array[14595]=30'd900139626;
array[14596]=30'd921150041;
array[14597]=30'd921150041;
array[14598]=30'd921150041;
array[14599]=30'd820526616;
array[14600]=30'd875034136;
array[14601]=30'd1033359876;
array[14602]=30'd1033359876;
array[14603]=30'd1033359876;
array[14604]=30'd1033359876;
array[14605]=30'd987238908;
array[14606]=30'd742923790;
array[14607]=30'd667440637;
array[14608]=30'd875034136;
array[14609]=30'd967280137;
array[14610]=30'd959928886;
array[14611]=30'd959928886;
array[14612]=30'd959928886;
array[14613]=30'd959928886;
array[14614]=30'd959928886;
array[14615]=30'd941029952;
array[14616]=30'd809995819;
array[14617]=30'd757545539;
array[14618]=30'd887567935;
array[14619]=30'd941029952;
array[14620]=30'd921150041;
array[14621]=30'd921150041;
array[14622]=30'd921150041;
array[14623]=30'd921150041;
array[14624]=30'd921150041;
array[14625]=30'd921150041;
array[14626]=30'd921150041;
array[14627]=30'd921150041;
array[14628]=30'd921150041;
array[14629]=30'd921150041;
array[14630]=30'd921150041;
array[14631]=30'd900139626;
array[14632]=30'd900139626;
array[14633]=30'd804758111;
array[14634]=30'd361192034;
array[14635]=30'd560346760;
array[14636]=30'd503733877;
array[14637]=30'd294104668;
array[14638]=30'd483946067;
array[14639]=30'd472478290;
array[14640]=30'd487155275;
array[14641]=30'd487155275;
array[14642]=30'd472478290;
array[14643]=30'd472478290;
array[14644]=30'd459884097;
array[14645]=30'd317277759;
array[14646]=30'd317277759;
array[14647]=30'd281613891;
array[14648]=30'd253299274;
array[14649]=30'd206107200;
array[14650]=30'd281613891;
array[14651]=30'd317277759;
array[14652]=30'd281613891;
array[14653]=30'd356077132;
array[14654]=30'd459884097;
array[14655]=30'd412701256;
array[14656]=30'd361277993;
array[14657]=30'd417793613;
array[14658]=30'd503733877;
array[14659]=30'd384241245;
array[14660]=30'd199687796;
array[14661]=30'd384241245;
array[14662]=30'd393770575;
array[14663]=30'd483946067;
array[14664]=30'd472478290;
array[14665]=30'd472478290;
array[14666]=30'd472478290;
array[14667]=30'd459884097;
array[14668]=30'd412701256;
array[14669]=30'd472478290;
array[14670]=30'd459884097;
array[14671]=30'd566784583;
array[14672]=30'd921150041;
array[14673]=30'd900139626;
array[14674]=30'd900139626;
array[14675]=30'd900139626;
array[14676]=30'd900139626;
array[14677]=30'd900139626;
array[14678]=30'd900139626;
array[14679]=30'd900139626;
array[14680]=30'd900139626;
array[14681]=30'd900139626;
array[14682]=30'd900139626;
array[14683]=30'd900139626;
array[14684]=30'd900139626;
array[14685]=30'd900139626;
array[14686]=30'd900139626;
array[14687]=30'd900139626;
array[14688]=30'd900139626;
array[14689]=30'd900139626;
array[14690]=30'd900139626;
array[14691]=30'd921150041;
array[14692]=30'd921150041;
array[14693]=30'd921150041;
array[14694]=30'd921150041;
array[14695]=30'd921150041;
array[14696]=30'd898098744;
array[14697]=30'd809995819;
array[14698]=30'd950544914;
array[14699]=30'd1033359876;
array[14700]=30'd1033359876;
array[14701]=30'd1004004888;
array[14702]=30'd910663171;
array[14703]=30'd742923790;
array[14704]=30'd985089582;
array[14705]=30'd959928886;
array[14706]=30'd959928886;
array[14707]=30'd959928886;
array[14708]=30'd959928886;
array[14709]=30'd959928886;
array[14710]=30'd959928886;
array[14711]=30'd959928886;
array[14712]=30'd959928886;
array[14713]=30'd916923947;
array[14714]=30'd757545539;
array[14715]=30'd941029952;
array[14716]=30'd921150041;
array[14717]=30'd921150041;
array[14718]=30'd921150041;
array[14719]=30'd921150041;
array[14720]=30'd921150041;
array[14721]=30'd921150041;
array[14722]=30'd921150041;
array[14723]=30'd921150041;
array[14724]=30'd921150041;
array[14725]=30'd921150041;
array[14726]=30'd900139626;
array[14727]=30'd900139626;
array[14728]=30'd900139626;
array[14729]=30'd549944915;
array[14730]=30'd451435107;
array[14731]=30'd453416554;
array[14732]=30'd503733877;
array[14733]=30'd352820791;
array[14734]=30'd518580800;
array[14735]=30'd472478290;
array[14736]=30'd487155275;
array[14737]=30'd487155275;
array[14738]=30'd487155275;
array[14739]=30'd472478290;
array[14740]=30'd472478290;
array[14741]=30'd472478290;
array[14742]=30'd459884097;
array[14743]=30'd459884097;
array[14744]=30'd412701256;
array[14745]=30'd281613891;
array[14746]=30'd459884097;
array[14747]=30'd459884097;
array[14748]=30'd459884097;
array[14749]=30'd412701256;
array[14750]=30'd412701256;
array[14751]=30'd356077132;
array[14752]=30'd431516230;
array[14753]=30'd482780758;
array[14754]=30'd453416554;
array[14755]=30'd294104668;
array[14756]=30'd245885528;
array[14757]=30'd361192034;
array[14758]=30'd451435107;
array[14759]=30'd459884097;
array[14760]=30'd472478290;
array[14761]=30'd472478290;
array[14762]=30'd459884097;
array[14763]=30'd412701256;
array[14764]=30'd472478290;
array[14765]=30'd472478290;
array[14766]=30'd472478290;
array[14767]=30'd412701256;
array[14768]=30'd840392271;
array[14769]=30'd921150041;
array[14770]=30'd900139626;
array[14771]=30'd900139626;
array[14772]=30'd900139626;
array[14773]=30'd900139626;
array[14774]=30'd900139626;
array[14775]=30'd900139626;
array[14776]=30'd900139626;
array[14777]=30'd900139626;
array[14778]=30'd900139626;
array[14779]=30'd900139626;
array[14780]=30'd900139626;
array[14781]=30'd900139626;
array[14782]=30'd900139626;
array[14783]=30'd900139626;
array[14784]=30'd900139626;
array[14785]=30'd900139626;
array[14786]=30'd900139626;
array[14787]=30'd921150041;
array[14788]=30'd921150041;
array[14789]=30'd921150041;
array[14790]=30'd921150041;
array[14791]=30'd921150041;
array[14792]=30'd921150041;
array[14793]=30'd921150041;
array[14794]=30'd809995819;
array[14795]=30'd809995819;
array[14796]=30'd967280137;
array[14797]=30'd935829023;
array[14798]=30'd679964212;
array[14799]=30'd898098744;
array[14800]=30'd985089582;
array[14801]=30'd959928886;
array[14802]=30'd959928886;
array[14803]=30'd959928886;
array[14804]=30'd959928886;
array[14805]=30'd959928886;
array[14806]=30'd959928886;
array[14807]=30'd959928886;
array[14808]=30'd959928886;
array[14809]=30'd959928886;
array[14810]=30'd757545539;
array[14811]=30'd887567935;
array[14812]=30'd921150041;
array[14813]=30'd921150041;
array[14814]=30'd921150041;
array[14815]=30'd921150041;
array[14816]=30'd921150041;
array[14817]=30'd921150041;
array[14818]=30'd921150041;
array[14819]=30'd921150041;
array[14820]=30'd900139626;
array[14821]=30'd900139626;
array[14822]=30'd921150041;
array[14823]=30'd921150041;
array[14824]=30'd804758111;
array[14825]=30'd431516230;
array[14826]=30'd483946067;
array[14827]=30'd393770575;
array[14828]=30'd451435107;
array[14829]=30'd339237463;
array[14830]=30'd483946067;
array[14831]=30'd472478290;
array[14832]=30'd487155275;
array[14833]=30'd487155275;
array[14834]=30'd487155275;
array[14835]=30'd487155275;
array[14836]=30'd472478290;
array[14837]=30'd472478290;
array[14838]=30'd472478290;
array[14839]=30'd472478290;
array[14840]=30'd459884097;
array[14841]=30'd412701256;
array[14842]=30'd472478290;
array[14843]=30'd472478290;
array[14844]=30'd472478290;
array[14845]=30'd472478290;
array[14846]=30'd472478290;
array[14847]=30'd459884097;
array[14848]=30'd459884097;
array[14849]=30'd393770575;
array[14850]=30'd453416554;
array[14851]=30'd294104668;
array[14852]=30'd393770575;
array[14853]=30'd302559805;
array[14854]=30'd431516230;
array[14855]=30'd472478290;
array[14856]=30'd472478290;
array[14857]=30'd472478290;
array[14858]=30'd412701256;
array[14859]=30'd459884097;
array[14860]=30'd472478290;
array[14861]=30'd472478290;
array[14862]=30'd472478290;
array[14863]=30'd459884097;
array[14864]=30'd698889775;
array[14865]=30'd921150041;
array[14866]=30'd900139626;
array[14867]=30'd900139626;
array[14868]=30'd900139626;
array[14869]=30'd900139626;
array[14870]=30'd900139626;
array[14871]=30'd900139626;
array[14872]=30'd900139626;
array[14873]=30'd921150041;
array[14874]=30'd921150041;
array[14875]=30'd921150041;
array[14876]=30'd921150041;
array[14877]=30'd921150041;
array[14878]=30'd921150041;
array[14879]=30'd921150041;
array[14880]=30'd921150041;
array[14881]=30'd900139626;
array[14882]=30'd921150041;
array[14883]=30'd921150041;
array[14884]=30'd921150041;
array[14885]=30'd921150041;
array[14886]=30'd921150041;
array[14887]=30'd921150041;
array[14888]=30'd921150041;
array[14889]=30'd921150041;
array[14890]=30'd921150041;
array[14891]=30'd898098744;
array[14892]=30'd778555959;
array[14893]=30'd679964212;
array[14894]=30'd617068069;
array[14895]=30'd959928886;
array[14896]=30'd959928886;
array[14897]=30'd959928886;
array[14898]=30'd959928886;
array[14899]=30'd959928886;
array[14900]=30'd959928886;
array[14901]=30'd959928886;
array[14902]=30'd959928886;
array[14903]=30'd959928886;
array[14904]=30'd959928886;
array[14905]=30'd959928886;
array[14906]=30'd809995819;
array[14907]=30'd887567935;
array[14908]=30'd921150041;
array[14909]=30'd921150041;
array[14910]=30'd921150041;
array[14911]=30'd921150041;
array[14912]=30'd921150041;
array[14913]=30'd921150041;
array[14914]=30'd921150041;
array[14915]=30'd921150041;
array[14916]=30'd921150041;
array[14917]=30'd921150041;
array[14918]=30'd921150041;
array[14919]=30'd887567935;
array[14920]=30'd506984008;
array[14921]=30'd472478290;
array[14922]=30'd472478290;
array[14923]=30'd483946067;
array[14924]=30'd339237463;
array[14925]=30'd339237463;
array[14926]=30'd393770575;
array[14927]=30'd459884097;
array[14928]=30'd487155275;
array[14929]=30'd487155275;
array[14930]=30'd487155275;
array[14931]=30'd487155275;
array[14932]=30'd487155275;
array[14933]=30'd472478290;
array[14934]=30'd472478290;
array[14935]=30'd472478290;
array[14936]=30'd412701256;
array[14937]=30'd472478290;
array[14938]=30'd472478290;
array[14939]=30'd472478290;
array[14940]=30'd472478290;
array[14941]=30'd472478290;
array[14942]=30'd472478290;
array[14943]=30'd472478290;
array[14944]=30'd459884097;
array[14945]=30'd339237463;
array[14946]=30'd339237463;
array[14947]=30'd393770575;
array[14948]=30'd483946067;
array[14949]=30'd361277993;
array[14950]=30'd356077132;
array[14951]=30'd472478290;
array[14952]=30'd472478290;
array[14953]=30'd459884097;
array[14954]=30'd412701256;
array[14955]=30'd472478290;
array[14956]=30'd472478290;
array[14957]=30'd459884097;
array[14958]=30'd472478290;
array[14959]=30'd459884097;
array[14960]=30'd566784583;
array[14961]=30'd921150041;
array[14962]=30'd900139626;
array[14963]=30'd900139626;
array[14964]=30'd900139626;
array[14965]=30'd900139626;
array[14966]=30'd921150041;
array[14967]=30'd900139626;
array[14968]=30'd921150041;
array[14969]=30'd921150041;
array[14970]=30'd935829023;
array[14971]=30'd935829023;
array[14972]=30'd875034136;
array[14973]=30'd855119352;
array[14974]=30'd855119352;
array[14975]=30'd875034136;
array[14976]=30'd921150041;
array[14977]=30'd921150041;
array[14978]=30'd921150041;
array[14979]=30'd921150041;
array[14980]=30'd921150041;
array[14981]=30'd921150041;
array[14982]=30'd921150041;
array[14983]=30'd921150041;
array[14984]=30'd921150041;
array[14985]=30'd921150041;
array[14986]=30'd921150041;
array[14987]=30'd921150041;
array[14988]=30'd921150041;
array[14989]=30'd921150041;
array[14990]=30'd679964212;
array[14991]=30'd959928886;
array[14992]=30'd959928886;
array[14993]=30'd959928886;
array[14994]=30'd959928886;
array[14995]=30'd959928886;
array[14996]=30'd959928886;
array[14997]=30'd959928886;
array[14998]=30'd959928886;
array[14999]=30'd959928886;
array[15000]=30'd959928886;
array[15001]=30'd959928886;
array[15002]=30'd809995819;
array[15003]=30'd757545539;
array[15004]=30'd887567935;
array[15005]=30'd921150041;
array[15006]=30'd921150041;
array[15007]=30'd921150041;
array[15008]=30'd921150041;
array[15009]=30'd921150041;
array[15010]=30'd921150041;
array[15011]=30'd921150041;
array[15012]=30'd921150041;
array[15013]=30'd921150041;
array[15014]=30'd898098744;
array[15015]=30'd506984008;
array[15016]=30'd483946067;
array[15017]=30'd472478290;
array[15018]=30'd487155275;
array[15019]=30'd487155275;
array[15020]=30'd393770575;
array[15021]=30'd302559805;
array[15022]=30'd431516230;
array[15023]=30'd472478290;
array[15024]=30'd472478290;
array[15025]=30'd487155275;
array[15026]=30'd487155275;
array[15027]=30'd487155275;
array[15028]=30'd487155275;
array[15029]=30'd472478290;
array[15030]=30'd472478290;
array[15031]=30'd459884097;
array[15032]=30'd412701256;
array[15033]=30'd472478290;
array[15034]=30'd472478290;
array[15035]=30'd472478290;
array[15036]=30'd472478290;
array[15037]=30'd472478290;
array[15038]=30'd472478290;
array[15039]=30'd472478290;
array[15040]=30'd472478290;
array[15041]=30'd356077132;
array[15042]=30'd302559805;
array[15043]=30'd483946067;
array[15044]=30'd472478290;
array[15045]=30'd459884097;
array[15046]=30'd317277759;
array[15047]=30'd459884097;
array[15048]=30'd472478290;
array[15049]=30'd412701256;
array[15050]=30'd472478290;
array[15051]=30'd472478290;
array[15052]=30'd472478290;
array[15053]=30'd472478290;
array[15054]=30'd472478290;
array[15055]=30'd472478290;
array[15056]=30'd483946067;
array[15057]=30'd921150041;
array[15058]=30'd921150041;
array[15059]=30'd921150041;
array[15060]=30'd921150041;
array[15061]=30'd921150041;
array[15062]=30'd921150041;
array[15063]=30'd921150041;
array[15064]=30'd1004004888;
array[15065]=30'd888658404;
array[15066]=30'd811098555;
array[15067]=30'd782796193;
array[15068]=30'd782796193;
array[15069]=30'd782796193;
array[15070]=30'd782796193;
array[15071]=30'd764964292;
array[15072]=30'd935829023;
array[15073]=30'd921150041;
array[15074]=30'd921150041;
array[15075]=30'd921150041;
array[15076]=30'd921150041;
array[15077]=30'd921150041;
array[15078]=30'd921150041;
array[15079]=30'd921150041;
array[15080]=30'd921150041;
array[15081]=30'd921150041;
array[15082]=30'd921150041;
array[15083]=30'd921150041;
array[15084]=30'd921150041;
array[15085]=30'd921150041;
array[15086]=30'd755499588;
array[15087]=30'd898098744;
array[15088]=30'd959928886;
array[15089]=30'd959928886;
array[15090]=30'd959928886;
array[15091]=30'd959928886;
array[15092]=30'd959928886;
array[15093]=30'd959928886;
array[15094]=30'd959928886;
array[15095]=30'd959928886;
array[15096]=30'd959928886;
array[15097]=30'd959928886;
array[15098]=30'd721911330;
array[15099]=30'd809995819;
array[15100]=30'd809995819;
array[15101]=30'd778555959;
array[15102]=30'd757545539;
array[15103]=30'd809995819;
array[15104]=30'd840392271;
array[15105]=30'd887567935;
array[15106]=30'd921150041;
array[15107]=30'd921150041;
array[15108]=30'd921150041;
array[15109]=30'd921150041;
array[15110]=30'd566784583;
array[15111]=30'd483946067;
array[15112]=30'd472478290;
array[15113]=30'd487155275;
array[15114]=30'd487155275;
array[15115]=30'd487155275;
array[15116]=30'd412701256;
array[15117]=30'd302559805;
array[15118]=30'd356077132;
array[15119]=30'd487155275;
array[15120]=30'd487155275;
array[15121]=30'd487155275;
array[15122]=30'd487155275;
array[15123]=30'd487155275;
array[15124]=30'd472478290;
array[15125]=30'd472478290;
array[15126]=30'd472478290;
array[15127]=30'd412701256;
array[15128]=30'd472478290;
array[15129]=30'd472478290;
array[15130]=30'd472478290;
array[15131]=30'd472478290;
array[15132]=30'd472478290;
array[15133]=30'd472478290;
array[15134]=30'd487155275;
array[15135]=30'd472478290;
array[15136]=30'd472478290;
array[15137]=30'd412701256;
array[15138]=30'd253299274;
array[15139]=30'd459884097;
array[15140]=30'd472478290;
array[15141]=30'd472478290;
array[15142]=30'd459884097;
array[15143]=30'd459884097;
array[15144]=30'd412701256;
array[15145]=30'd412701256;
array[15146]=30'd472478290;
array[15147]=30'd472478290;
array[15148]=30'd472478290;
array[15149]=30'd459884097;
array[15150]=30'd472478290;
array[15151]=30'd472478290;
array[15152]=30'd412701256;
array[15153]=30'd840392271;
array[15154]=30'd921150041;
array[15155]=30'd921150041;
array[15156]=30'd921150041;
array[15157]=30'd921150041;
array[15158]=30'd921150041;
array[15159]=30'd1004004888;
array[15160]=30'd926429685;
array[15161]=30'd764964292;
array[15162]=30'd811098555;
array[15163]=30'd849905057;
array[15164]=30'd849905057;
array[15165]=30'd906527146;
array[15166]=30'd945318330;
array[15167]=30'd811098555;
array[15168]=30'd888658404;
array[15169]=30'd935829023;
array[15170]=30'd941029952;
array[15171]=30'd941029952;
array[15172]=30'd921150041;
array[15173]=30'd921150041;
array[15174]=30'd921150041;
array[15175]=30'd921150041;
array[15176]=30'd921150041;
array[15177]=30'd921150041;
array[15178]=30'd921150041;
array[15179]=30'd921150041;
array[15180]=30'd921150041;
array[15181]=30'd921150041;
array[15182]=30'd921150041;
array[15183]=30'd778555959;
array[15184]=30'd840392271;
array[15185]=30'd959928886;
array[15186]=30'd959928886;
array[15187]=30'd959928886;
array[15188]=30'd959928886;
array[15189]=30'd959928886;
array[15190]=30'd959928886;
array[15191]=30'd959928886;
array[15192]=30'd959928886;
array[15193]=30'd916923947;
array[15194]=30'd778555959;
array[15195]=30'd1004004888;
array[15196]=30'd1033359876;
array[15197]=30'd1033359876;
array[15198]=30'd1004004888;
array[15199]=30'd967280137;
array[15200]=30'd875034136;
array[15201]=30'd809995819;
array[15202]=30'd778555959;
array[15203]=30'd757545539;
array[15204]=30'd757545539;
array[15205]=30'd583554612;
array[15206]=30'd453527098;
array[15207]=30'd487155275;
array[15208]=30'd487155275;
array[15209]=30'd472478290;
array[15210]=30'd472478290;
array[15211]=30'd459884097;
array[15212]=30'd412701256;
array[15213]=30'd472478290;
array[15214]=30'd356077132;
array[15215]=30'd459884097;
array[15216]=30'd472478290;
array[15217]=30'd487155275;
array[15218]=30'd487155275;
array[15219]=30'd472478290;
array[15220]=30'd472478290;
array[15221]=30'd472478290;
array[15222]=30'd459884097;
array[15223]=30'd412701256;
array[15224]=30'd472478290;
array[15225]=30'd472478290;
array[15226]=30'd472478290;
array[15227]=30'd472478290;
array[15228]=30'd472478290;
array[15229]=30'd472478290;
array[15230]=30'd487155275;
array[15231]=30'd472478290;
array[15232]=30'd459884097;
array[15233]=30'd483946067;
array[15234]=30'd302559805;
array[15235]=30'd483946067;
array[15236]=30'd487155275;
array[15237]=30'd472478290;
array[15238]=30'd472478290;
array[15239]=30'd472478290;
array[15240]=30'd356077132;
array[15241]=30'd472478290;
array[15242]=30'd472478290;
array[15243]=30'd472478290;
array[15244]=30'd472478290;
array[15245]=30'd472478290;
array[15246]=30'd472478290;
array[15247]=30'd472478290;
array[15248]=30'd459884097;
array[15249]=30'd733487691;
array[15250]=30'd921150041;
array[15251]=30'd921150041;
array[15252]=30'd921150041;
array[15253]=30'd921150041;
array[15254]=30'd959928886;
array[15255]=30'd950544914;
array[15256]=30'd811098555;
array[15257]=30'd833137031;
array[15258]=30'd943234452;
array[15259]=30'd849905057;
array[15260]=30'd782796193;
array[15261]=30'd869807552;
array[15262]=30'd1000883648;
array[15263]=30'd906527146;
array[15264]=30'd811098555;
array[15265]=30'd888658404;
array[15266]=30'd935829023;
array[15267]=30'd941029952;
array[15268]=30'd941029952;
array[15269]=30'd921150041;
array[15270]=30'd921150041;
array[15271]=30'd921150041;
array[15272]=30'd921150041;
array[15273]=30'd921150041;
array[15274]=30'd921150041;
array[15275]=30'd921150041;
array[15276]=30'd921150041;
array[15277]=30'd921150041;
array[15278]=30'd921150041;
array[15279]=30'd921150041;
array[15280]=30'd840392271;
array[15281]=30'd757545539;
array[15282]=30'd862402083;
array[15283]=30'd935829023;
array[15284]=30'd809995819;
array[15285]=30'd809995819;
array[15286]=30'd916923947;
array[15287]=30'd959928886;
array[15288]=30'd959928886;
array[15289]=30'd721911330;
array[15290]=30'd679964212;
array[15291]=30'd844591615;
array[15292]=30'd967280137;
array[15293]=30'd1004004888;
array[15294]=30'd1033359876;
array[15295]=30'd1033359876;
array[15296]=30'd1033359876;
array[15297]=30'd1033359876;
array[15298]=30'd1033359876;
array[15299]=30'd1004004888;
array[15300]=30'd950544914;
array[15301]=30'd624454176;
array[15302]=30'd400051721;
array[15303]=30'd414764563;
array[15304]=30'd414764563;
array[15305]=30'd481862174;
array[15306]=30'd412701256;
array[15307]=30'd412701256;
array[15308]=30'd496575016;
array[15309]=30'd472478290;
array[15310]=30'd472478290;
array[15311]=30'd459884097;
array[15312]=30'd472478290;
array[15313]=30'd487155275;
array[15314]=30'd472478290;
array[15315]=30'd472478290;
array[15316]=30'd472478290;
array[15317]=30'd472478290;
array[15318]=30'd356077132;
array[15319]=30'd459884097;
array[15320]=30'd472478290;
array[15321]=30'd472478290;
array[15322]=30'd472478290;
array[15323]=30'd472478290;
array[15324]=30'd472478290;
array[15325]=30'd472478290;
array[15326]=30'd487155275;
array[15327]=30'd472478290;
array[15328]=30'd542677555;
array[15329]=30'd840392271;
array[15330]=30'd642228804;
array[15331]=30'd655912516;
array[15332]=30'd459884097;
array[15333]=30'd472478290;
array[15334]=30'd472478290;
array[15335]=30'd459884097;
array[15336]=30'd317277759;
array[15337]=30'd459884097;
array[15338]=30'd412701256;
array[15339]=30'd459884097;
array[15340]=30'd472478290;
array[15341]=30'd472478290;
array[15342]=30'd472478290;
array[15343]=30'd472478290;
array[15344]=30'd472478290;
array[15345]=30'd542677555;
array[15346]=30'd921150041;
array[15347]=30'd921150041;
array[15348]=30'd921150041;
array[15349]=30'd959928886;
array[15350]=30'd1004004888;
array[15351]=30'd832058842;
array[15352]=30'd768126344;
array[15353]=30'd885566856;
array[15354]=30'd833137031;
array[15355]=30'd768126344;
array[15356]=30'd768126344;
array[15357]=30'd782796193;
array[15358]=30'd945318330;
array[15359]=30'd945318330;
array[15360]=30'd906527146;
array[15361]=30'd832058842;
array[15362]=30'd946320871;
array[15363]=30'd935829023;
array[15364]=30'd916923947;
array[15365]=30'd921150041;
array[15366]=30'd921150041;
array[15367]=30'd921150041;
array[15368]=30'd921150041;
array[15369]=30'd921150041;
array[15370]=30'd921150041;
array[15371]=30'd921150041;
array[15372]=30'd921150041;
array[15373]=30'd921150041;
array[15374]=30'd921150041;
array[15375]=30'd921150041;
array[15376]=30'd921150041;
array[15377]=30'd921150041;
array[15378]=30'd804758111;
array[15379]=30'd595020337;
array[15380]=30'd887567935;
array[15381]=30'd935829023;
array[15382]=30'd809995819;
array[15383]=30'd721911330;
array[15384]=30'd778555959;
array[15385]=30'd862402083;
array[15386]=30'd935829023;
array[15387]=30'd721911330;
array[15388]=30'd651672075;
array[15389]=30'd721911330;
array[15390]=30'd721911330;
array[15391]=30'd778555959;
array[15392]=30'd809995819;
array[15393]=30'd935829023;
array[15394]=30'd1004004888;
array[15395]=30'd1033359876;
array[15396]=30'd1033359876;
array[15397]=30'd708323812;
array[15398]=30'd491266512;
array[15399]=30'd491266512;
array[15400]=30'd491266512;
array[15401]=30'd443016687;
array[15402]=30'd372793832;
array[15403]=30'd361277993;
array[15404]=30'd412701256;
array[15405]=30'd459884097;
array[15406]=30'd487155275;
array[15407]=30'd472478290;
array[15408]=30'd472478290;
array[15409]=30'd472478290;
array[15410]=30'd487155275;
array[15411]=30'd472478290;
array[15412]=30'd356077132;
array[15413]=30'd412701256;
array[15414]=30'd412701256;
array[15415]=30'd472478290;
array[15416]=30'd472478290;
array[15417]=30'd487155275;
array[15418]=30'd472478290;
array[15419]=30'd472478290;
array[15420]=30'd487155275;
array[15421]=30'd472478290;
array[15422]=30'd472478290;
array[15423]=30'd518580800;
array[15424]=30'd840392271;
array[15425]=30'd642228804;
array[15426]=30'd713478705;
array[15427]=30'd642228804;
array[15428]=30'd483946067;
array[15429]=30'd459884097;
array[15430]=30'd496575016;
array[15431]=30'd412701256;
array[15432]=30'd820526616;
array[15433]=30'd935829023;
array[15434]=30'd898098744;
array[15435]=30'd542677555;
array[15436]=30'd459884097;
array[15437]=30'd472478290;
array[15438]=30'd472478290;
array[15439]=30'd472478290;
array[15440]=30'd472478290;
array[15441]=30'd459884097;
array[15442]=30'd733487691;
array[15443]=30'd959928886;
array[15444]=30'd959928886;
array[15445]=30'd1004004888;
array[15446]=30'd926429685;
array[15447]=30'd764964292;
array[15448]=30'd833137031;
array[15449]=30'd768126344;
array[15450]=30'd768126344;
array[15451]=30'd849905057;
array[15452]=30'd906527146;
array[15453]=30'd849905057;
array[15454]=30'd945318330;
array[15455]=30'd849905057;
array[15456]=30'd869807552;
array[15457]=30'd832058842;
array[15458]=30'd964180446;
array[15459]=30'd888658404;
array[15460]=30'd910663171;
array[15461]=30'd916923947;
array[15462]=30'd921150041;
array[15463]=30'd921150041;
array[15464]=30'd921150041;
array[15465]=30'd921150041;
array[15466]=30'd921150041;
array[15467]=30'd921150041;
array[15468]=30'd921150041;
array[15469]=30'd921150041;
array[15470]=30'd921150041;
array[15471]=30'd921150041;
array[15472]=30'd921150041;
array[15473]=30'd921150041;
array[15474]=30'd921150041;
array[15475]=30'd809995819;
array[15476]=30'd809995819;
array[15477]=30'd959928886;
array[15478]=30'd959928886;
array[15479]=30'd862402083;
array[15480]=30'd757545539;
array[15481]=30'd985089582;
array[15482]=30'd959928886;
array[15483]=30'd959928886;
array[15484]=30'd757545539;
array[15485]=30'd887567935;
array[15486]=30'd959928886;
array[15487]=30'd921150041;
array[15488]=30'd898098744;
array[15489]=30'd809995819;
array[15490]=30'd506984008;
array[15491]=30'd583554612;
array[15492]=30'd667440637;
array[15493]=30'd531143170;
array[15494]=30'd457732594;
array[15495]=30'd491266512;
array[15496]=30'd491266512;
array[15497]=30'd477614540;
array[15498]=30'd477614540;
array[15499]=30'd491266512;
array[15500]=30'd443016687;
array[15501]=30'd400051721;
array[15502]=30'd414764563;
array[15503]=30'd481862174;
array[15504]=30'd459884097;
array[15505]=30'd459884097;
array[15506]=30'd472478290;
array[15507]=30'd472478290;
array[15508]=30'd412701256;
array[15509]=30'd356077132;
array[15510]=30'd459884097;
array[15511]=30'd472478290;
array[15512]=30'd472478290;
array[15513]=30'd472478290;
array[15514]=30'd487155275;
array[15515]=30'd472478290;
array[15516]=30'd472478290;
array[15517]=30'd487155275;
array[15518]=30'd487155275;
array[15519]=30'd518580800;
array[15520]=30'd733487691;
array[15521]=30'd757545539;
array[15522]=30'd794232376;
array[15523]=30'd721911330;
array[15524]=30'd481862174;
array[15525]=30'd481862174;
array[15526]=30'd481862174;
array[15527]=30'd414764563;
array[15528]=30'd809995819;
array[15529]=30'd809995819;
array[15530]=30'd809995819;
array[15531]=30'd583554612;
array[15532]=30'd481862174;
array[15533]=30'd459884097;
array[15534]=30'd472478290;
array[15535]=30'd472478290;
array[15536]=30'd472478290;
array[15537]=30'd459884097;
array[15538]=30'd412701256;
array[15539]=30'd857219651;
array[15540]=30'd959928886;
array[15541]=30'd1004004888;
array[15542]=30'd855119352;
array[15543]=30'd782796193;
array[15544]=30'd885566856;
array[15545]=30'd768126344;
array[15546]=30'd782796193;
array[15547]=30'd906527146;
array[15548]=30'd979923369;
array[15549]=30'd945318330;
array[15550]=30'd849905057;
array[15551]=30'd782796193;
array[15552]=30'd855016073;
array[15553]=30'd855016073;
array[15554]=30'd855016073;
array[15555]=30'd855016073;
array[15556]=30'd855016073;
array[15557]=30'd855016073;
array[15558]=30'd855016073;
array[15559]=30'd855016073;
array[15560]=30'd855016073;
array[15561]=30'd855016073;
array[15562]=30'd855016073;
array[15563]=30'd855016073;
array[15564]=30'd855016073;
array[15565]=30'd855016073;
array[15566]=30'd855016073;
array[15567]=30'd855016073;
array[15568]=30'd855016073;
array[15569]=30'd855016073;
array[15570]=30'd855016073;
array[15571]=30'd855016073;
array[15572]=30'd855016073;
array[15573]=30'd855016073;
array[15574]=30'd855016073;
array[15575]=30'd855016073;
array[15576]=30'd855016073;
array[15577]=30'd855016073;
array[15578]=30'd855016073;
array[15579]=30'd855016073;
array[15580]=30'd855016073;
array[15581]=30'd879170165;
array[15582]=30'd883367490;
array[15583]=30'd824630873;
array[15584]=30'd824630873;
array[15585]=30'd855016073;
array[15586]=30'd855016073;
array[15587]=30'd855016073;
array[15588]=30'd855016073;
array[15589]=30'd855016073;
array[15590]=30'd855016073;
array[15591]=30'd855016073;
array[15592]=30'd855016073;
array[15593]=30'd855016073;
array[15594]=30'd855016073;
array[15595]=30'd730239616;
array[15596]=30'd463850128;
array[15597]=30'd463850128;
array[15598]=30'd556097214;
array[15599]=30'd601183923;
array[15600]=30'd601183923;
array[15601]=30'd539297481;
array[15602]=30'd633679565;
array[15603]=30'd633679565;
array[15604]=30'd601183923;
array[15605]=30'd601183923;
array[15606]=30'd630512344;
array[15607]=30'd630512344;
array[15608]=30'd601183923;
array[15609]=30'd651585154;
array[15610]=30'd523632283;
array[15611]=30'd601183923;
array[15612]=30'd630512344;
array[15613]=30'd630512344;
array[15614]=30'd630512344;
array[15615]=30'd630512344;
array[15616]=30'd630512344;
array[15617]=30'd630512344;
array[15618]=30'd646252225;
array[15619]=30'd630512344;
array[15620]=30'd630512344;
array[15621]=30'd601183923;
array[15622]=30'd394645149;
array[15623]=30'd601183923;
array[15624]=30'd646252225;
array[15625]=30'd633679565;
array[15626]=30'd630512344;
array[15627]=30'd630512344;
array[15628]=30'd630512344;
array[15629]=30'd630512344;
array[15630]=30'd601183923;
array[15631]=30'd583395966;
array[15632]=30'd883367490;
array[15633]=30'd883367490;
array[15634]=30'd824630873;
array[15635]=30'd816210575;
array[15636]=30'd816210575;
array[15637]=30'd816210575;
array[15638]=30'd855016073;
array[15639]=30'd816210575;
array[15640]=30'd855016073;
array[15641]=30'd855016073;
array[15642]=30'd855016073;
array[15643]=30'd855016073;
array[15644]=30'd855016073;
array[15645]=30'd855016073;
array[15646]=30'd855016073;
array[15647]=30'd879170165;
array[15648]=30'd855016073;
array[15649]=30'd855016073;
array[15650]=30'd855016073;
array[15651]=30'd855016073;
array[15652]=30'd855016073;
array[15653]=30'd855016073;
array[15654]=30'd855016073;
array[15655]=30'd855016073;
array[15656]=30'd855016073;
array[15657]=30'd855016073;
array[15658]=30'd855016073;
array[15659]=30'd855016073;
array[15660]=30'd855016073;
array[15661]=30'd855016073;
array[15662]=30'd855016073;
array[15663]=30'd855016073;
array[15664]=30'd855016073;
array[15665]=30'd855016073;
array[15666]=30'd855016073;
array[15667]=30'd855016073;
array[15668]=30'd855016073;
array[15669]=30'd855016073;
array[15670]=30'd855016073;
array[15671]=30'd855016073;
array[15672]=30'd855016073;
array[15673]=30'd855016073;
array[15674]=30'd855016073;
array[15675]=30'd855016073;
array[15676]=30'd855016073;
array[15677]=30'd855016073;
array[15678]=30'd855016073;
array[15679]=30'd855016073;
array[15680]=30'd855016073;
array[15681]=30'd855016073;
array[15682]=30'd855016073;
array[15683]=30'd855016073;
array[15684]=30'd855016073;
array[15685]=30'd855016073;
array[15686]=30'd855016073;
array[15687]=30'd855016073;
array[15688]=30'd855016073;
array[15689]=30'd855016073;
array[15690]=30'd816210575;
array[15691]=30'd583395966;
array[15692]=30'd452327079;
array[15693]=30'd611709603;
array[15694]=30'd444947126;
array[15695]=30'd601183923;
array[15696]=30'd518350503;
array[15697]=30'd601183923;
array[15698]=30'd646252225;
array[15699]=30'd646252225;
array[15700]=30'd486895284;
array[15701]=30'd646252225;
array[15702]=30'd630512344;
array[15703]=30'd646252225;
array[15704]=30'd548775573;
array[15705]=30'd794239590;
array[15706]=30'd527849061;
array[15707]=30'd637892242;
array[15708]=30'd630512344;
array[15709]=30'd630512344;
array[15710]=30'd630512344;
array[15711]=30'd630512344;
array[15712]=30'd630512344;
array[15713]=30'd630512344;
array[15714]=30'd633679565;
array[15715]=30'd630512344;
array[15716]=30'd630512344;
array[15717]=30'd633679565;
array[15718]=30'd394645149;
array[15719]=30'd497425057;
array[15720]=30'd646252225;
array[15721]=30'd633679565;
array[15722]=30'd630512344;
array[15723]=30'd630512344;
array[15724]=30'd633679565;
array[15725]=30'd633679565;
array[15726]=30'd646252225;
array[15727]=30'd611709603;
array[15728]=30'd665233987;
array[15729]=30'd824630873;
array[15730]=30'd824630873;
array[15731]=30'd816210575;
array[15732]=30'd816210575;
array[15733]=30'd855016073;
array[15734]=30'd816210575;
array[15735]=30'd855016073;
array[15736]=30'd855016073;
array[15737]=30'd855016073;
array[15738]=30'd855016073;
array[15739]=30'd855016073;
array[15740]=30'd879170165;
array[15741]=30'd879170165;
array[15742]=30'd900141674;
array[15743]=30'd959930934;
array[15744]=30'd816210575;
array[15745]=30'd855016073;
array[15746]=30'd855016073;
array[15747]=30'd855016073;
array[15748]=30'd855016073;
array[15749]=30'd855016073;
array[15750]=30'd855016073;
array[15751]=30'd855016073;
array[15752]=30'd855016073;
array[15753]=30'd855016073;
array[15754]=30'd855016073;
array[15755]=30'd855016073;
array[15756]=30'd855016073;
array[15757]=30'd855016073;
array[15758]=30'd855016073;
array[15759]=30'd855016073;
array[15760]=30'd855016073;
array[15761]=30'd855016073;
array[15762]=30'd855016073;
array[15763]=30'd855016073;
array[15764]=30'd855016073;
array[15765]=30'd855016073;
array[15766]=30'd855016073;
array[15767]=30'd855016073;
array[15768]=30'd855016073;
array[15769]=30'd855016073;
array[15770]=30'd855016073;
array[15771]=30'd855016073;
array[15772]=30'd855016073;
array[15773]=30'd855016073;
array[15774]=30'd855016073;
array[15775]=30'd855016073;
array[15776]=30'd855016073;
array[15777]=30'd855016073;
array[15778]=30'd855016073;
array[15779]=30'd855016073;
array[15780]=30'd855016073;
array[15781]=30'd855016073;
array[15782]=30'd855016073;
array[15783]=30'd855016073;
array[15784]=30'd855016073;
array[15785]=30'd855016073;
array[15786]=30'd779516542;
array[15787]=30'd452327079;
array[15788]=30'd463850128;
array[15789]=30'd601183923;
array[15790]=30'd486895284;
array[15791]=30'd646252225;
array[15792]=30'd486895284;
array[15793]=30'd646252225;
array[15794]=30'd646252225;
array[15795]=30'd601183923;
array[15796]=30'd486895284;
array[15797]=30'd646252225;
array[15798]=30'd630512344;
array[15799]=30'd556097214;
array[15800]=30'd730239616;
array[15801]=30'd824630873;
array[15802]=30'd527849061;
array[15803]=30'd668323493;
array[15804]=30'd633679565;
array[15805]=30'd630512344;
array[15806]=30'd630512344;
array[15807]=30'd630512344;
array[15808]=30'd630512344;
array[15809]=30'd630512344;
array[15810]=30'd646252225;
array[15811]=30'd630512344;
array[15812]=30'd630512344;
array[15813]=30'd633679565;
array[15814]=30'd518350503;
array[15815]=30'd354789034;
array[15816]=30'd601183923;
array[15817]=30'd633679565;
array[15818]=30'd630512344;
array[15819]=30'd630512344;
array[15820]=30'd539297481;
array[15821]=30'd601183923;
array[15822]=30'd646252225;
array[15823]=30'd601183923;
array[15824]=30'd523632283;
array[15825]=30'd824630873;
array[15826]=30'd824630873;
array[15827]=30'd855016073;
array[15828]=30'd855016073;
array[15829]=30'd855016073;
array[15830]=30'd816210575;
array[15831]=30'd816210575;
array[15832]=30'd855016073;
array[15833]=30'd855016073;
array[15834]=30'd855016073;
array[15835]=30'd879170165;
array[15836]=30'd922198619;
array[15837]=30'd979844654;
array[15838]=30'd936883742;
array[15839]=30'd872938009;
array[15840]=30'd855016073;
array[15841]=30'd855016073;
array[15842]=30'd855016073;
array[15843]=30'd855016073;
array[15844]=30'd855016073;
array[15845]=30'd855016073;
array[15846]=30'd855016073;
array[15847]=30'd855016073;
array[15848]=30'd855016073;
array[15849]=30'd855016073;
array[15850]=30'd855016073;
array[15851]=30'd855016073;
array[15852]=30'd855016073;
array[15853]=30'd855016073;
array[15854]=30'd879170165;
array[15855]=30'd879170165;
array[15856]=30'd879170165;
array[15857]=30'd883367490;
array[15858]=30'd883367490;
array[15859]=30'd824630873;
array[15860]=30'd879170165;
array[15861]=30'd879170165;
array[15862]=30'd879170165;
array[15863]=30'd855016073;
array[15864]=30'd855016073;
array[15865]=30'd855016073;
array[15866]=30'd855016073;
array[15867]=30'd855016073;
array[15868]=30'd855016073;
array[15869]=30'd855016073;
array[15870]=30'd855016073;
array[15871]=30'd855016073;
array[15872]=30'd855016073;
array[15873]=30'd855016073;
array[15874]=30'd855016073;
array[15875]=30'd855016073;
array[15876]=30'd855016073;
array[15877]=30'd855016073;
array[15878]=30'd855016073;
array[15879]=30'd855016073;
array[15880]=30'd855016073;
array[15881]=30'd855016073;
array[15882]=30'd651585154;
array[15883]=30'd463850128;
array[15884]=30'd583395966;
array[15885]=30'd556097214;
array[15886]=30'd556097214;
array[15887]=30'd601183923;
array[15888]=30'd518350503;
array[15889]=30'd646252225;
array[15890]=30'd646252225;
array[15891]=30'd486895284;
array[15892]=30'd556097214;
array[15893]=30'd646252225;
array[15894]=30'd646252225;
array[15895]=30'd583395966;
array[15896]=30'd941029952;
array[15897]=30'd824630873;
array[15898]=30'd557205073;
array[15899]=30'd637892242;
array[15900]=30'd601183923;
array[15901]=30'd646252225;
array[15902]=30'd630512344;
array[15903]=30'd633679565;
array[15904]=30'd556097214;
array[15905]=30'd630512344;
array[15906]=30'd630512344;
array[15907]=30'd630512344;
array[15908]=30'd630512344;
array[15909]=30'd633679565;
array[15910]=30'd556097214;
array[15911]=30'd289797789;
array[15912]=30'd611709603;
array[15913]=30'd646252225;
array[15914]=30'd630512344;
array[15915]=30'd630512344;
array[15916]=30'd630512344;
array[15917]=30'd518350503;
array[15918]=30'd646252225;
array[15919]=30'd646252225;
array[15920]=30'd548775573;
array[15921]=30'd779516542;
array[15922]=30'd816210575;
array[15923]=30'd855016073;
array[15924]=30'd855016073;
array[15925]=30'd855016073;
array[15926]=30'd855016073;
array[15927]=30'd855016073;
array[15928]=30'd855016073;
array[15929]=30'd855016073;
array[15930]=30'd855016073;
array[15931]=30'd879170165;
array[15932]=30'd898098744;
array[15933]=30'd820526616;
array[15934]=30'd777516526;
array[15935]=30'd777516526;
array[15936]=30'd855016073;
array[15937]=30'd855016073;
array[15938]=30'd855016073;
array[15939]=30'd855016073;
array[15940]=30'd855016073;
array[15941]=30'd855016073;
array[15942]=30'd855016073;
array[15943]=30'd855016073;
array[15944]=30'd855016073;
array[15945]=30'd855016073;
array[15946]=30'd855016073;
array[15947]=30'd879170165;
array[15948]=30'd900141674;
array[15949]=30'd959930934;
array[15950]=30'd936883742;
array[15951]=30'd872938009;
array[15952]=30'd855121400;
array[15953]=30'd871846383;
array[15954]=30'd839346691;
array[15955]=30'd804744750;
array[15956]=30'd859252262;
array[15957]=30'd916919852;
array[15958]=30'd916919852;
array[15959]=30'd804744750;
array[15960]=30'd842497613;
array[15961]=30'd855016073;
array[15962]=30'd855016073;
array[15963]=30'd855016073;
array[15964]=30'd855016073;
array[15965]=30'd855016073;
array[15966]=30'd855016073;
array[15967]=30'd855016073;
array[15968]=30'd855016073;
array[15969]=30'd855016073;
array[15970]=30'd855016073;
array[15971]=30'd855016073;
array[15972]=30'd855016073;
array[15973]=30'd855016073;
array[15974]=30'd855016073;
array[15975]=30'd855016073;
array[15976]=30'd855016073;
array[15977]=30'd816210575;
array[15978]=30'd497425057;
array[15979]=30'd463850128;
array[15980]=30'd637892242;
array[15981]=30'd486895284;
array[15982]=30'd601183923;
array[15983]=30'd548775573;
array[15984]=30'd556097214;
array[15985]=30'd633679565;
array[15986]=30'd646252225;
array[15987]=30'd497425057;
array[15988]=30'd556097214;
array[15989]=30'd646252225;
array[15990]=30'd601183923;
array[15991]=30'd751243845;
array[15992]=30'd941029952;
array[15993]=30'd883367490;
array[15994]=30'd527849061;
array[15995]=30'd637892242;
array[15996]=30'd444947126;
array[15997]=30'd637892242;
array[15998]=30'd646252225;
array[15999]=30'd646252225;
array[16000]=30'd427157133;
array[16001]=30'd646252225;
array[16002]=30'd630512344;
array[16003]=30'd630512344;
array[16004]=30'd630512344;
array[16005]=30'd601183923;
array[16006]=30'd601183923;
array[16007]=30'd322308749;
array[16008]=30'd523632283;
array[16009]=30'd646252225;
array[16010]=30'd633679565;
array[16011]=30'd630512344;
array[16012]=30'd630512344;
array[16013]=30'd539297481;
array[16014]=30'd646252225;
array[16015]=30'd646252225;
array[16016]=30'd601183923;
array[16017]=30'd695644807;
array[16018]=30'd855016073;
array[16019]=30'd855016073;
array[16020]=30'd855016073;
array[16021]=30'd855016073;
array[16022]=30'd855016073;
array[16023]=30'd855016073;
array[16024]=30'd855016073;
array[16025]=30'd855016073;
array[16026]=30'd855016073;
array[16027]=30'd879170165;
array[16028]=30'd842497613;
array[16029]=30'd804744750;
array[16030]=30'd839346691;
array[16031]=30'd859252262;
array[16032]=30'd855016073;
array[16033]=30'd855016073;
array[16034]=30'd855016073;
array[16035]=30'd855016073;
array[16036]=30'd855016073;
array[16037]=30'd855016073;
array[16038]=30'd855016073;
array[16039]=30'd855016073;
array[16040]=30'd855016073;
array[16041]=30'd879170165;
array[16042]=30'd879170165;
array[16043]=30'd900141674;
array[16044]=30'd959930934;
array[16045]=30'd916977147;
array[16046]=30'd809003452;
array[16047]=30'd767069629;
array[16048]=30'd741905818;
array[16049]=30'd741905818;
array[16050]=30'd589828536;
array[16051]=30'd414702010;
array[16052]=30'd422024669;
array[16053]=30'd694663659;
array[16054]=30'd916977147;
array[16055]=30'd777516526;
array[16056]=30'd839346691;
array[16057]=30'd883367490;
array[16058]=30'd855016073;
array[16059]=30'd855016073;
array[16060]=30'd855016073;
array[16061]=30'd855016073;
array[16062]=30'd855016073;
array[16063]=30'd855016073;
array[16064]=30'd855016073;
array[16065]=30'd855016073;
array[16066]=30'd855016073;
array[16067]=30'd855016073;
array[16068]=30'd855016073;
array[16069]=30'd855016073;
array[16070]=30'd855016073;
array[16071]=30'd855016073;
array[16072]=30'd855016073;
array[16073]=30'd730239616;
array[16074]=30'd503735925;
array[16075]=30'd463850128;
array[16076]=30'd668323493;
array[16077]=30'd444947126;
array[16078]=30'd668323493;
array[16079]=30'd518350503;
array[16080]=30'd601183923;
array[16081]=30'd646252225;
array[16082]=30'd556097214;
array[16083]=30'd583395966;
array[16084]=30'd611709603;
array[16085]=30'd668323493;
array[16086]=30'd548775573;
array[16087]=30'd883367490;
array[16088]=30'd941029952;
array[16089]=30'd883367490;
array[16090]=30'd510044739;
array[16091]=30'd614845038;
array[16092]=30'd614845038;
array[16093]=30'd559303301;
array[16094]=30'd646252225;
array[16095]=30'd646252225;
array[16096]=30'd497425057;
array[16097]=30'd548775573;
array[16098]=30'd646252225;
array[16099]=30'd630512344;
array[16100]=30'd630512344;
array[16101]=30'd486895284;
array[16102]=30'd601183923;
array[16103]=30'd322308749;
array[16104]=30'd463850128;
array[16105]=30'd646252225;
array[16106]=30'd630512344;
array[16107]=30'd630512344;
array[16108]=30'd630512344;
array[16109]=30'd601183923;
array[16110]=30'd556097214;
array[16111]=30'd646252225;
array[16112]=30'd646252225;
array[16113]=30'd583395966;
array[16114]=30'd855016073;
array[16115]=30'd855016073;
array[16116]=30'd855016073;
array[16117]=30'd855016073;
array[16118]=30'd855016073;
array[16119]=30'd855016073;
array[16120]=30'd855016073;
array[16121]=30'd855016073;
array[16122]=30'd855016073;
array[16123]=30'd855016073;
array[16124]=30'd855016073;
array[16125]=30'd879170165;
array[16126]=30'd879170165;
array[16127]=30'd900141674;
array[16128]=30'd855016073;
array[16129]=30'd855016073;
array[16130]=30'd855016073;
array[16131]=30'd855016073;
array[16132]=30'd855016073;
array[16133]=30'd855016073;
array[16134]=30'd855016073;
array[16135]=30'd855016073;
array[16136]=30'd855016073;
array[16137]=30'd879170165;
array[16138]=30'd900141674;
array[16139]=30'd959930934;
array[16140]=30'd916977147;
array[16141]=30'd767069629;
array[16142]=30'd849905057;
array[16143]=30'd908629408;
array[16144]=30'd792242589;
array[16145]=30'd661135811;
array[16146]=30'd414702010;
array[16147]=30'd461875644;
array[16148]=30'd422024669;
array[16149]=30'd422024669;
array[16150]=30'd737670674;
array[16151]=30'd661135811;
array[16152]=30'd735537629;
array[16153]=30'd859252262;
array[16154]=30'd855016073;
array[16155]=30'd855016073;
array[16156]=30'd855016073;
array[16157]=30'd855016073;
array[16158]=30'd855016073;
array[16159]=30'd855016073;
array[16160]=30'd855016073;
array[16161]=30'd855016073;
array[16162]=30'd855016073;
array[16163]=30'd855016073;
array[16164]=30'd855016073;
array[16165]=30'd855016073;
array[16166]=30'd855016073;
array[16167]=30'd855016073;
array[16168]=30'd855016073;
array[16169]=30'd651585154;
array[16170]=30'd548775573;
array[16171]=30'd523632283;
array[16172]=30'd668323493;
array[16173]=30'd444947126;
array[16174]=30'd668323493;
array[16175]=30'd463850128;
array[16176]=30'd668323493;
array[16177]=30'd601183923;
array[16178]=30'd559303301;
array[16179]=30'd695644807;
array[16180]=30'd583395966;
array[16181]=30'd601183923;
array[16182]=30'd624350812;
array[16183]=30'd941029952;
array[16184]=30'd941029952;
array[16185]=30'd916919852;
array[16186]=30'd539404850;
array[16187]=30'd614845038;
array[16188]=30'd751243845;
array[16189]=30'd527849061;
array[16190]=30'd637892242;
array[16191]=30'd668323493;
array[16192]=30'd651585154;
array[16193]=30'd568787568;
array[16194]=30'd637892242;
array[16195]=30'd646252225;
array[16196]=30'd633679565;
array[16197]=30'd444947126;
array[16198]=30'd556097214;
array[16199]=30'd362168943;
array[16200]=30'd373711515;
array[16201]=30'd637892242;
array[16202]=30'd633679565;
array[16203]=30'd630512344;
array[16204]=30'd630512344;
array[16205]=30'd633679565;
array[16206]=30'd518350503;
array[16207]=30'd646252225;
array[16208]=30'd646252225;
array[16209]=30'd548775573;
array[16210]=30'd816210575;
array[16211]=30'd855016073;
array[16212]=30'd855016073;
array[16213]=30'd855016073;
array[16214]=30'd855016073;
array[16215]=30'd855016073;
array[16216]=30'd855016073;
array[16217]=30'd855016073;
array[16218]=30'd855016073;
array[16219]=30'd855016073;
array[16220]=30'd855016073;
array[16221]=30'd855016073;
array[16222]=30'd855016073;
array[16223]=30'd922198619;
array[16224]=30'd855016073;
array[16225]=30'd855016073;
array[16226]=30'd855016073;
array[16227]=30'd855016073;
array[16228]=30'd855016073;
array[16229]=30'd855016073;
array[16230]=30'd855016073;
array[16231]=30'd879170165;
array[16232]=30'd879170165;
array[16233]=30'd900141674;
array[16234]=30'd959930934;
array[16235]=30'd916977147;
array[16236]=30'd809003452;
array[16237]=30'd829990281;
array[16238]=30'd876132737;
array[16239]=30'd741905818;
array[16240]=30'd553137612;
array[16241]=30'd323471799;
array[16242]=30'd323471799;
array[16243]=30'd323471799;
array[16244]=30'd279425485;
array[16245]=30'd241691107;
array[16246]=30'd279425485;
array[16247]=30'd323471799;
array[16248]=30'd422024669;
array[16249]=30'd761730564;
array[16250]=30'd824630873;
array[16251]=30'd855016073;
array[16252]=30'd855016073;
array[16253]=30'd855016073;
array[16254]=30'd855016073;
array[16255]=30'd855016073;
array[16256]=30'd855016073;
array[16257]=30'd855016073;
array[16258]=30'd855016073;
array[16259]=30'd855016073;
array[16260]=30'd855016073;
array[16261]=30'd855016073;
array[16262]=30'd855016073;
array[16263]=30'd855016073;
array[16264]=30'd855016073;
array[16265]=30'd559303301;
array[16266]=30'd548775573;
array[16267]=30'd548775573;
array[16268]=30'd668323493;
array[16269]=30'd444947126;
array[16270]=30'd601183923;
array[16271]=30'd373711515;
array[16272]=30'd637892242;
array[16273]=30'd611709603;
array[16274]=30'd624350812;
array[16275]=30'd792119862;
array[16276]=30'd583395966;
array[16277]=30'd611709603;
array[16278]=30'd751243845;
array[16279]=30'd959930934;
array[16280]=30'd959930934;
array[16281]=30'd941029952;
array[16282]=30'd624350812;
array[16283]=30'd568787568;
array[16284]=30'd824630873;
array[16285]=30'd751243845;
array[16286]=30'd583395966;
array[16287]=30'd668323493;
array[16288]=30'd559303301;
array[16289]=30'd792119862;
array[16290]=30'd583395966;
array[16291]=30'd637892242;
array[16292]=30'd646252225;
array[16293]=30'd518350503;
array[16294]=30'd497425057;
array[16295]=30'd427157133;
array[16296]=30'd362168943;
array[16297]=30'd637892242;
array[16298]=30'd633679565;
array[16299]=30'd630512344;
array[16300]=30'd630512344;
array[16301]=30'd633679565;
array[16302]=30'd518350503;
array[16303]=30'd633679565;
array[16304]=30'd646252225;
array[16305]=30'd518350503;
array[16306]=30'd816210575;
array[16307]=30'd855016073;
array[16308]=30'd855016073;
array[16309]=30'd855016073;
array[16310]=30'd855016073;
array[16311]=30'd855016073;
array[16312]=30'd855016073;
array[16313]=30'd855016073;
array[16314]=30'd855016073;
array[16315]=30'd855016073;
array[16316]=30'd855016073;
array[16317]=30'd855016073;
array[16318]=30'd879170165;
array[16319]=30'd883367490;
array[16320]=30'd855016073;
array[16321]=30'd855016073;
array[16322]=30'd855016073;
array[16323]=30'd855016073;
array[16324]=30'd855016073;
array[16325]=30'd855016073;
array[16326]=30'd879170165;
array[16327]=30'd879170165;
array[16328]=30'd879170165;
array[16329]=30'd922198619;
array[16330]=30'd936883742;
array[16331]=30'd767069629;
array[16332]=30'd829990281;
array[16333]=30'd792242589;
array[16334]=30'd766030218;
array[16335]=30'd792242589;
array[16336]=30'd753420739;
array[16337]=30'd414702010;
array[16338]=30'd461875644;
array[16339]=30'd461875644;
array[16340]=30'd359126474;
array[16341]=30'd359126474;
array[16342]=30'd461875644;
array[16343]=30'd461875644;
array[16344]=30'd422024669;
array[16345]=30'd722945572;
array[16346]=30'd665233987;
array[16347]=30'd651585154;
array[16348]=30'd695644807;
array[16349]=30'd779516542;
array[16350]=30'd855016073;
array[16351]=30'd855016073;
array[16352]=30'd855016073;
array[16353]=30'd855016073;
array[16354]=30'd855016073;
array[16355]=30'd855016073;
array[16356]=30'd855016073;
array[16357]=30'd855016073;
array[16358]=30'd855016073;
array[16359]=30'd855016073;
array[16360]=30'd816210575;
array[16361]=30'd497425057;
array[16362]=30'd548775573;
array[16363]=30'd548775573;
array[16364]=30'd601183923;
array[16365]=30'd373711515;
array[16366]=30'd583395966;
array[16367]=30'd433488509;
array[16368]=30'd614845038;
array[16369]=30'd611709603;
array[16370]=30'd751243845;
array[16371]=30'd824630873;
array[16372]=30'd503735925;
array[16373]=30'd583395966;
array[16374]=30'd824630873;
array[16375]=30'd959930934;
array[16376]=30'd959930934;
array[16377]=30'd959930934;
array[16378]=30'd792119862;
array[16379]=30'd527849061;
array[16380]=30'd792119862;
array[16381]=30'd916919852;
array[16382]=30'd527849061;
array[16383]=30'd637892242;
array[16384]=30'd503735925;
array[16385]=30'd883367490;
array[16386]=30'd557205073;
array[16387]=30'd637892242;
array[16388]=30'd601183923;
array[16389]=30'd583395966;
array[16390]=30'd503735925;
array[16391]=30'd568787568;
array[16392]=30'd484882002;
array[16393]=30'd637892242;
array[16394]=30'd633679565;
array[16395]=30'd633679565;
array[16396]=30'd630512344;
array[16397]=30'd633679565;
array[16398]=30'd539297481;
array[16399]=30'd633679565;
array[16400]=30'd646252225;
array[16401]=30'd556097214;
array[16402]=30'd779516542;
array[16403]=30'd855016073;
array[16404]=30'd855016073;
array[16405]=30'd816210575;
array[16406]=30'd855016073;
array[16407]=30'd855016073;
array[16408]=30'd855016073;
array[16409]=30'd855016073;
array[16410]=30'd855016073;
array[16411]=30'd855016073;
array[16412]=30'd855016073;
array[16413]=30'd855016073;
array[16414]=30'd855016073;
array[16415]=30'd855016073;
array[16416]=30'd855016073;
array[16417]=30'd855016073;
array[16418]=30'd855016073;
array[16419]=30'd855016073;
array[16420]=30'd855016073;
array[16421]=30'd855016073;
array[16422]=30'd879170165;
array[16423]=30'd879170165;
array[16424]=30'd879170165;
array[16425]=30'd959930934;
array[16426]=30'd855121400;
array[16427]=30'd809003452;
array[16428]=30'd876132737;
array[16429]=30'd766030218;
array[16430]=30'd809003452;
array[16431]=30'd893925805;
array[16432]=30'd871910847;
array[16433]=30'd414702010;
array[16434]=30'd479712691;
array[16435]=30'd461875644;
array[16436]=30'd359126474;
array[16437]=30'd359126474;
array[16438]=30'd479712691;
array[16439]=30'd461875644;
array[16440]=30'd492300766;
array[16441]=30'd859252262;
array[16442]=30'd824630873;
array[16443]=30'd855016073;
array[16444]=30'd816210575;
array[16445]=30'd730239616;
array[16446]=30'd681987696;
array[16447]=30'd695644807;
array[16448]=30'd816210575;
array[16449]=30'd855016073;
array[16450]=30'd855016073;
array[16451]=30'd855016073;
array[16452]=30'd855016073;
array[16453]=30'd855016073;
array[16454]=30'd855016073;
array[16455]=30'd855016073;
array[16456]=30'd779516542;
array[16457]=30'd548775573;
array[16458]=30'd556097214;
array[16459]=30'd518350503;
array[16460]=30'd611709603;
array[16461]=30'd322308749;
array[16462]=30'd503735925;
array[16463]=30'd665233987;
array[16464]=30'd557205073;
array[16465]=30'd527849061;
array[16466]=30'd665233987;
array[16467]=30'd804744750;
array[16468]=30'd510044739;
array[16469]=30'd503735925;
array[16470]=30'd794239590;
array[16471]=30'd959930934;
array[16472]=30'd959930934;
array[16473]=30'd959930934;
array[16474]=30'd883367490;
array[16475]=30'd484882002;
array[16476]=30'd679961142;
array[16477]=30'd679961142;
array[16478]=30'd708220465;
array[16479]=30'd559303301;
array[16480]=30'd503735925;
array[16481]=30'd665233987;
array[16482]=30'd624350812;
array[16483]=30'd583395966;
array[16484]=30'd637892242;
array[16485]=30'd593953387;
array[16486]=30'd568787568;
array[16487]=30'd571952708;
array[16488]=30'd665233987;
array[16489]=30'd614845038;
array[16490]=30'd646252225;
array[16491]=30'd601183923;
array[16492]=30'd633679565;
array[16493]=30'd633679565;
array[16494]=30'd556097214;
array[16495]=30'd601183923;
array[16496]=30'd646252225;
array[16497]=30'd556097214;
array[16498]=30'd779516542;
array[16499]=30'd855016073;
array[16500]=30'd855016073;
array[16501]=30'd855016073;
array[16502]=30'd855016073;
array[16503]=30'd855016073;
array[16504]=30'd855016073;
array[16505]=30'd855016073;
array[16506]=30'd855016073;
array[16507]=30'd855016073;
array[16508]=30'd855016073;
array[16509]=30'd855016073;
array[16510]=30'd855016073;
array[16511]=30'd855016073;
array[16512]=30'd855016073;
array[16513]=30'd855016073;
array[16514]=30'd855016073;
array[16515]=30'd855016073;
array[16516]=30'd855016073;
array[16517]=30'd855016073;
array[16518]=30'd879170165;
array[16519]=30'd879170165;
array[16520]=30'd879170165;
array[16521]=30'd959930934;
array[16522]=30'd855121400;
array[16523]=30'd809003452;
array[16524]=30'd908629408;
array[16525]=30'd792242589;
array[16526]=30'd809003452;
array[16527]=30'd945318330;
array[16528]=30'd809003452;
array[16529]=30'd394764738;
array[16530]=30'd479712691;
array[16531]=30'd448250284;
array[16532]=30'd394764738;
array[16533]=30'd372750770;
array[16534]=30'd461875644;
array[16535]=30'd461875644;
array[16536]=30'd684132856;
array[16537]=30'd842497613;
array[16538]=30'd855016073;
array[16539]=30'd855016073;
array[16540]=30'd855016073;
array[16541]=30'd855016073;
array[16542]=30'd855016073;
array[16543]=30'd816210575;
array[16544]=30'd730239616;
array[16545]=30'd695644807;
array[16546]=30'd779516542;
array[16547]=30'd855016073;
array[16548]=30'd855016073;
array[16549]=30'd855016073;
array[16550]=30'd855016073;
array[16551]=30'd855016073;
array[16552]=30'd695644807;
array[16553]=30'd583395966;
array[16554]=30'd601183923;
array[16555]=30'd518350503;
array[16556]=30'd556097214;
array[16557]=30'd477520516;
array[16558]=30'd484882002;
array[16559]=30'd792119862;
array[16560]=30'd484882002;
array[16561]=30'd557205073;
array[16562]=30'd941029952;
array[16563]=30'd941029952;
array[16564]=30'd679961142;
array[16565]=30'd548890196;
array[16566]=30'd941029952;
array[16567]=30'd959930934;
array[16568]=30'd959930934;
array[16569]=30'd959930934;
array[16570]=30'd941029952;
array[16571]=30'd751243845;
array[16572]=30'd679961142;
array[16573]=30'd959930934;
array[16574]=30'd941029952;
array[16575]=30'd665233987;
array[16576]=30'd527849061;
array[16577]=30'd916919852;
array[16578]=30'd859252262;
array[16579]=30'd527849061;
array[16580]=30'd614845038;
array[16581]=30'd679961142;
array[16582]=30'd641176139;
array[16583]=30'd679961142;
array[16584]=30'd792119862;
array[16585]=30'd583395966;
array[16586]=30'd601183923;
array[16587]=30'd601183923;
array[16588]=30'd633679565;
array[16589]=30'd633679565;
array[16590]=30'd601183923;
array[16591]=30'd556097214;
array[16592]=30'd633679565;
array[16593]=30'd601183923;
array[16594]=30'd730239616;
array[16595]=30'd855016073;
array[16596]=30'd855016073;
array[16597]=30'd855016073;
array[16598]=30'd855016073;
array[16599]=30'd855016073;
array[16600]=30'd855016073;
array[16601]=30'd855016073;
array[16602]=30'd855016073;
array[16603]=30'd855016073;
array[16604]=30'd855016073;
array[16605]=30'd855016073;
array[16606]=30'd855016073;
array[16607]=30'd855016073;
array[16608]=30'd855016073;
array[16609]=30'd855016073;
array[16610]=30'd855016073;
array[16611]=30'd855016073;
array[16612]=30'd855016073;
array[16613]=30'd855016073;
array[16614]=30'd879170165;
array[16615]=30'd879170165;
array[16616]=30'd879170165;
array[16617]=30'd922198619;
array[16618]=30'd872938009;
array[16619]=30'd753420739;
array[16620]=30'd871910847;
array[16621]=30'd871910847;
array[16622]=30'd778590630;
array[16623]=30'd778590630;
array[16624]=30'd661135811;
array[16625]=30'd414702010;
array[16626]=30'd479712691;
array[16627]=30'd479712691;
array[16628]=30'd461875644;
array[16629]=30'd448250284;
array[16630]=30'd461875644;
array[16631]=30'd422024669;
array[16632]=30'd792119862;
array[16633]=30'd824630873;
array[16634]=30'd855016073;
array[16635]=30'd855016073;
array[16636]=30'd855016073;
array[16637]=30'd855016073;
array[16638]=30'd855016073;
array[16639]=30'd855016073;
array[16640]=30'd855016073;
array[16641]=30'd855016073;
array[16642]=30'd779516542;
array[16643]=30'd695644807;
array[16644]=30'd779516542;
array[16645]=30'd855016073;
array[16646]=30'd855016073;
array[16647]=30'd855016073;
array[16648]=30'd651585154;
array[16649]=30'd637892242;
array[16650]=30'd646252225;
array[16651]=30'd452327079;
array[16652]=30'd548775573;
array[16653]=30'd707208791;
array[16654]=30'd417795660;
array[16655]=30'd679961142;
array[16656]=30'd583428668;
array[16657]=30'd548890196;
array[16658]=30'd959930934;
array[16659]=30'd959930934;
array[16660]=30'd883367490;
array[16661]=30'd571952708;
array[16662]=30'd959930934;
array[16663]=30'd959930934;
array[16664]=30'd959930934;
array[16665]=30'd959930934;
array[16666]=30'd941029952;
array[16667]=30'd941029952;
array[16668]=30'd768057919;
array[16669]=30'd959930934;
array[16670]=30'd959930934;
array[16671]=30'd883367490;
array[16672]=30'd539404850;
array[16673]=30'd916919852;
array[16674]=30'd959930934;
array[16675]=30'd751243845;
array[16676]=30'd484882002;
array[16677]=30'd751243845;
array[16678]=30'd722945572;
array[16679]=30'd768057919;
array[16680]=30'd751243845;
array[16681]=30'd484882002;
array[16682]=30'd637892242;
array[16683]=30'd556097214;
array[16684]=30'd601183923;
array[16685]=30'd633679565;
array[16686]=30'd601183923;
array[16687]=30'd539297481;
array[16688]=30'd633679565;
array[16689]=30'd601183923;
array[16690]=30'd730239616;
array[16691]=30'd855016073;
array[16692]=30'd855016073;
array[16693]=30'd855016073;
array[16694]=30'd855016073;
array[16695]=30'd855016073;
array[16696]=30'd855016073;
array[16697]=30'd855016073;
array[16698]=30'd855016073;
array[16699]=30'd855016073;
array[16700]=30'd855016073;
array[16701]=30'd855016073;
array[16702]=30'd855016073;
array[16703]=30'd855016073;
array[16704]=30'd855016073;
array[16705]=30'd855016073;
array[16706]=30'd855016073;
array[16707]=30'd855016073;
array[16708]=30'd855016073;
array[16709]=30'd855016073;
array[16710]=30'd879170165;
array[16711]=30'd879170165;
array[16712]=30'd879170165;
array[16713]=30'd900141674;
array[16714]=30'd936883742;
array[16715]=30'd767069629;
array[16716]=30'd792195525;
array[16717]=30'd894969309;
array[16718]=30'd815247846;
array[16719]=30'd777516526;
array[16720]=30'd619182551;
array[16721]=30'd414702010;
array[16722]=30'd479712691;
array[16723]=30'd479712691;
array[16724]=30'd479712691;
array[16725]=30'd414702010;
array[16726]=30'd394764738;
array[16727]=30'd422024669;
array[16728]=30'd859252262;
array[16729]=30'd824630873;
array[16730]=30'd855016073;
array[16731]=30'd855016073;
array[16732]=30'd879170165;
array[16733]=30'd794239590;
array[16734]=30'd593953387;
array[16735]=30'd730239616;
array[16736]=30'd855016073;
array[16737]=30'd855016073;
array[16738]=30'd855016073;
array[16739]=30'd855016073;
array[16740]=30'd779516542;
array[16741]=30'd695644807;
array[16742]=30'd779516542;
array[16743]=30'd855016073;
array[16744]=30'd559303301;
array[16745]=30'd637892242;
array[16746]=30'd646252225;
array[16747]=30'd518350503;
array[16748]=30'd523632283;
array[16749]=30'd751243845;
array[16750]=30'd468145703;
array[16751]=30'd941029952;
array[16752]=30'd883367490;
array[16753]=30'd571952708;
array[16754]=30'd959930934;
array[16755]=30'd959930934;
array[16756]=30'd959930934;
array[16757]=30'd916919852;
array[16758]=30'd959930934;
array[16759]=30'd959930934;
array[16760]=30'd959930934;
array[16761]=30'd959930934;
array[16762]=30'd979844654;
array[16763]=30'd959930934;
array[16764]=30'd959930934;
array[16765]=30'd959930934;
array[16766]=30'd959930934;
array[16767]=30'd959930934;
array[16768]=30'd883367490;
array[16769]=30'd941029952;
array[16770]=30'd959930934;
array[16771]=30'd883367490;
array[16772]=30'd510044739;
array[16773]=30'd859252262;
array[16774]=30'd597116464;
array[16775]=30'd804744750;
array[16776]=30'd442989058;
array[16777]=30'd491162135;
array[16778]=30'd457612903;
array[16779]=30'd523632283;
array[16780]=30'd601183923;
array[16781]=30'd633679565;
array[16782]=30'd633679565;
array[16783]=30'd556097214;
array[16784]=30'd633679565;
array[16785]=30'd601183923;
array[16786]=30'd730239616;
array[16787]=30'd855016073;
array[16788]=30'd855016073;
array[16789]=30'd855016073;
array[16790]=30'd855016073;
array[16791]=30'd855016073;
array[16792]=30'd855016073;
array[16793]=30'd855016073;
array[16794]=30'd855016073;
array[16795]=30'd855016073;
array[16796]=30'd855016073;
array[16797]=30'd855016073;
array[16798]=30'd855016073;
array[16799]=30'd855016073;
array[16800]=30'd855016073;
array[16801]=30'd855016073;
array[16802]=30'd855016073;
array[16803]=30'd855016073;
array[16804]=30'd855016073;
array[16805]=30'd879170165;
array[16806]=30'd855016073;
array[16807]=30'd879170165;
array[16808]=30'd879170165;
array[16809]=30'd879170165;
array[16810]=30'd959930934;
array[16811]=30'd855121400;
array[16812]=30'd753420739;
array[16813]=30'd832062938;
array[16814]=30'd894969309;
array[16815]=30'd855121400;
array[16816]=30'd586684918;
array[16817]=30'd461875644;
array[16818]=30'd479712691;
array[16819]=30'd490193319;
array[16820]=30'd479712691;
array[16821]=30'd461875644;
array[16822]=30'd394764738;
array[16823]=30'd504834577;
array[16824]=30'd635883032;
array[16825]=30'd681987696;
array[16826]=30'd779516542;
array[16827]=30'd824630873;
array[16828]=30'd571952708;
array[16829]=30'd396849695;
array[16830]=30'd468145703;
array[16831]=30'd597116464;
array[16832]=30'd883367490;
array[16833]=30'd855016073;
array[16834]=30'd855016073;
array[16835]=30'd855016073;
array[16836]=30'd855016073;
array[16837]=30'd855016073;
array[16838]=30'd779516542;
array[16839]=30'd651585154;
array[16840]=30'd457612903;
array[16841]=30'd668323493;
array[16842]=30'd646252225;
array[16843]=30'd601183923;
array[16844]=30'd427157133;
array[16845]=30'd751243845;
array[16846]=30'd883367490;
array[16847]=30'd959930934;
array[16848]=30'd959930934;
array[16849]=30'd883367490;
array[16850]=30'd959930934;
array[16851]=30'd959930934;
array[16852]=30'd959930934;
array[16853]=30'd959930934;
array[16854]=30'd959930934;
array[16855]=30'd959930934;
array[16856]=30'd959930934;
array[16857]=30'd959930934;
array[16858]=30'd979844654;
array[16859]=30'd979844654;
array[16860]=30'd959930934;
array[16861]=30'd959930934;
array[16862]=30'd959930934;
array[16863]=30'd959930934;
array[16864]=30'd959930934;
array[16865]=30'd979844654;
array[16866]=30'd959930934;
array[16867]=30'd959930934;
array[16868]=30'd916919852;
array[16869]=30'd959930934;
array[16870]=30'd859252262;
array[16871]=30'd804744750;
array[16872]=30'd650619404;
array[16873]=30'd815247846;
array[16874]=30'd449215039;
array[16875]=30'd484816502;
array[16876]=30'd601183923;
array[16877]=30'd633679565;
array[16878]=30'd633679565;
array[16879]=30'd556097214;
array[16880]=30'd630512344;
array[16881]=30'd556097214;
array[16882]=30'd779516542;
array[16883]=30'd855016073;
array[16884]=30'd855016073;
array[16885]=30'd855016073;
array[16886]=30'd855016073;
array[16887]=30'd855016073;
array[16888]=30'd855016073;
array[16889]=30'd855016073;
array[16890]=30'd855016073;
array[16891]=30'd855016073;
array[16892]=30'd855016073;
array[16893]=30'd855016073;
array[16894]=30'd855016073;
array[16895]=30'd855016073;
array[16896]=30'd855016073;
array[16897]=30'd855016073;
array[16898]=30'd855016073;
array[16899]=30'd855016073;
array[16900]=30'd855016073;
array[16901]=30'd855016073;
array[16902]=30'd879170165;
array[16903]=30'd879170165;
array[16904]=30'd879170165;
array[16905]=30'd879170165;
array[16906]=30'd898098744;
array[16907]=30'd898098744;
array[16908]=30'd785935846;
array[16909]=30'd809003452;
array[16910]=30'd832062938;
array[16911]=30'd832062938;
array[16912]=30'd553137612;
array[16913]=30'd461875644;
array[16914]=30'd479712691;
array[16915]=30'd490193319;
array[16916]=30'd479712691;
array[16917]=30'd461875644;
array[16918]=30'd422024669;
array[16919]=30'd792119862;
array[16920]=30'd842497613;
array[16921]=30'd794239590;
array[16922]=30'd527922743;
array[16923]=30'd333946399;
array[16924]=30'd371683842;
array[16925]=30'd422024669;
array[16926]=30'd475492838;
array[16927]=30'd597116464;
array[16928]=30'd883367490;
array[16929]=30'd855016073;
array[16930]=30'd855016073;
array[16931]=30'd855016073;
array[16932]=30'd855016073;
array[16933]=30'd855016073;
array[16934]=30'd855016073;
array[16935]=30'd816210575;
array[16936]=30'd457612903;
array[16937]=30'd548775573;
array[16938]=30'd601183923;
array[16939]=30'd601183923;
array[16940]=30'd548775573;
array[16941]=30'd768057919;
array[16942]=30'd959930934;
array[16943]=30'd959930934;
array[16944]=30'd959930934;
array[16945]=30'd959930934;
array[16946]=30'd883367490;
array[16947]=30'd883367490;
array[16948]=30'd883367490;
array[16949]=30'd959930934;
array[16950]=30'd959930934;
array[16951]=30'd959930934;
array[16952]=30'd959930934;
array[16953]=30'd959930934;
array[16954]=30'd959930934;
array[16955]=30'd959930934;
array[16956]=30'd959930934;
array[16957]=30'd959930934;
array[16958]=30'd959930934;
array[16959]=30'd959930934;
array[16960]=30'd959930934;
array[16961]=30'd959930934;
array[16962]=30'd959930934;
array[16963]=30'd959930934;
array[16964]=30'd959930934;
array[16965]=30'd959930934;
array[16966]=30'd959930934;
array[16967]=30'd872938009;
array[16968]=30'd650619404;
array[16969]=30'd777516526;
array[16970]=30'd510044739;
array[16971]=30'd484816502;
array[16972]=30'd637892242;
array[16973]=30'd646252225;
array[16974]=30'd633679565;
array[16975]=30'd556097214;
array[16976]=30'd630512344;
array[16977]=30'd556097214;
array[16978]=30'd779516542;
array[16979]=30'd855016073;
array[16980]=30'd855016073;
array[16981]=30'd855016073;
array[16982]=30'd855016073;
array[16983]=30'd855016073;
array[16984]=30'd855016073;
array[16985]=30'd855016073;
array[16986]=30'd855016073;
array[16987]=30'd855016073;
array[16988]=30'd855016073;
array[16989]=30'd855016073;
array[16990]=30'd855016073;
array[16991]=30'd855016073;
array[16992]=30'd855016073;
array[16993]=30'd855016073;
array[16994]=30'd855016073;
array[16995]=30'd855016073;
array[16996]=30'd879170165;
array[16997]=30'd855016073;
array[16998]=30'd879170165;
array[16999]=30'd879170165;
array[17000]=30'd879170165;
array[17001]=30'd879170165;
array[17002]=30'd879170165;
array[17003]=30'd898098744;
array[17004]=30'd872938009;
array[17005]=30'd785935846;
array[17006]=30'd792195525;
array[17007]=30'd753420739;
array[17008]=30'd461875644;
array[17009]=30'd461875644;
array[17010]=30'd479712691;
array[17011]=30'd490193319;
array[17012]=30'd479712691;
array[17013]=30'd448250284;
array[17014]=30'd504834577;
array[17015]=30'd883367490;
array[17016]=30'd824630873;
array[17017]=30'd679961142;
array[17018]=30'd442989058;
array[17019]=30'd475492838;
array[17020]=30'd414702010;
array[17021]=30'd359126474;
array[17022]=30'd279425485;
array[17023]=30'd665233987;
array[17024]=30'd824630873;
array[17025]=30'd855016073;
array[17026]=30'd855016073;
array[17027]=30'd855016073;
array[17028]=30'd855016073;
array[17029]=30'd855016073;
array[17030]=30'd855016073;
array[17031]=30'd855016073;
array[17032]=30'd559303301;
array[17033]=30'd548775573;
array[17034]=30'd486895284;
array[17035]=30'd486895284;
array[17036]=30'd611709603;
array[17037]=30'd751243845;
array[17038]=30'd959930934;
array[17039]=30'd959930934;
array[17040]=30'd859252262;
array[17041]=30'd722945572;
array[17042]=30'd722945572;
array[17043]=30'd859252262;
array[17044]=30'd804744750;
array[17045]=30'd804744750;
array[17046]=30'd959930934;
array[17047]=30'd979844654;
array[17048]=30'd979844654;
array[17049]=30'd959930934;
array[17050]=30'd959930934;
array[17051]=30'd959930934;
array[17052]=30'd959930934;
array[17053]=30'd916919852;
array[17054]=30'd804744750;
array[17055]=30'd722945572;
array[17056]=30'd722945572;
array[17057]=30'd768057919;
array[17058]=30'd916919852;
array[17059]=30'd959930934;
array[17060]=30'd959930934;
array[17061]=30'd959930934;
array[17062]=30'd959930934;
array[17063]=30'd859252262;
array[17064]=30'd468145703;
array[17065]=30'd504834577;
array[17066]=30'd557205073;
array[17067]=30'd484816502;
array[17068]=30'd601183923;
array[17069]=30'd646252225;
array[17070]=30'd633679565;
array[17071]=30'd556097214;
array[17072]=30'd633679565;
array[17073]=30'd518350503;
array[17074]=30'd816210575;
array[17075]=30'd855016073;
array[17076]=30'd855016073;
array[17077]=30'd855016073;
array[17078]=30'd855016073;
array[17079]=30'd855016073;
array[17080]=30'd855016073;
array[17081]=30'd855016073;
array[17082]=30'd855016073;
array[17083]=30'd855016073;
array[17084]=30'd855016073;
array[17085]=30'd855016073;
array[17086]=30'd855016073;
array[17087]=30'd855016073;
array[17088]=30'd855016073;
array[17089]=30'd855016073;
array[17090]=30'd855016073;
array[17091]=30'd855016073;
array[17092]=30'd879170165;
array[17093]=30'd879170165;
array[17094]=30'd879170165;
array[17095]=30'd879170165;
array[17096]=30'd879170165;
array[17097]=30'd879170165;
array[17098]=30'd900141674;
array[17099]=30'd959930934;
array[17100]=30'd916977147;
array[17101]=30'd815247846;
array[17102]=30'd871846383;
array[17103]=30'd839346691;
array[17104]=30'd441989592;
array[17105]=30'd479712691;
array[17106]=30'd479712691;
array[17107]=30'd490193319;
array[17108]=30'd479712691;
array[17109]=30'd448250284;
array[17110]=30'd650619404;
array[17111]=30'd883367490;
array[17112]=30'd679961142;
array[17113]=30'd442989058;
array[17114]=30'd492300766;
array[17115]=30'd479712691;
array[17116]=30'd448250284;
array[17117]=30'd394764738;
array[17118]=30'd442989058;
array[17119]=30'd751243845;
array[17120]=30'd681987696;
array[17121]=30'd816210575;
array[17122]=30'd855016073;
array[17123]=30'd855016073;
array[17124]=30'd855016073;
array[17125]=30'd855016073;
array[17126]=30'd855016073;
array[17127]=30'd855016073;
array[17128]=30'd559303301;
array[17129]=30'd637892242;
array[17130]=30'd601183923;
array[17131]=30'd419779260;
array[17132]=30'd637892242;
array[17133]=30'd624350812;
array[17134]=30'd941029952;
array[17135]=30'd768057919;
array[17136]=30'd768057919;
array[17137]=30'd737670674;
array[17138]=30'd468145703;
array[17139]=30'd333946399;
array[17140]=30'd597116464;
array[17141]=30'd916919852;
array[17142]=30'd959930934;
array[17143]=30'd979844654;
array[17144]=30'd979844654;
array[17145]=30'd959930934;
array[17146]=30'd959930934;
array[17147]=30'd959930934;
array[17148]=30'd941029952;
array[17149]=30'd751243845;
array[17150]=30'd804744750;
array[17151]=30'd722945572;
array[17152]=30'd679961142;
array[17153]=30'd722945572;
array[17154]=30'd679961142;
array[17155]=30'd722945572;
array[17156]=30'd916919852;
array[17157]=30'd959930934;
array[17158]=30'd959930934;
array[17159]=30'd936883742;
array[17160]=30'd722945572;
array[17161]=30'd527849061;
array[17162]=30'd614845038;
array[17163]=30'd452327079;
array[17164]=30'd646252225;
array[17165]=30'd646252225;
array[17166]=30'd601183923;
array[17167]=30'd556097214;
array[17168]=30'd646252225;
array[17169]=30'd548775573;
array[17170]=30'd855016073;
array[17171]=30'd855016073;
array[17172]=30'd855016073;
array[17173]=30'd855016073;
array[17174]=30'd855016073;
array[17175]=30'd855016073;
array[17176]=30'd855016073;
array[17177]=30'd855016073;
array[17178]=30'd855016073;
array[17179]=30'd855016073;
array[17180]=30'd855016073;
array[17181]=30'd855016073;
array[17182]=30'd855016073;
array[17183]=30'd855016073;
array[17184]=30'd855016073;
array[17185]=30'd855016073;
array[17186]=30'd855016073;
array[17187]=30'd855016073;
array[17188]=30'd879170165;
array[17189]=30'd879170165;
array[17190]=30'd879170165;
array[17191]=30'd879170165;
array[17192]=30'd879170165;
array[17193]=30'd900141674;
array[17194]=30'd959930934;
array[17195]=30'd996656669;
array[17196]=30'd832062938;
array[17197]=30'd815247846;
array[17198]=30'd936883742;
array[17199]=30'd916977147;
array[17200]=30'd422024669;
array[17201]=30'd479712691;
array[17202]=30'd490193319;
array[17203]=30'd490193319;
array[17204]=30'd490193319;
array[17205]=30'd414702010;
array[17206]=30'd761730564;
array[17207]=30'd613923367;
array[17208]=30'd442989058;
array[17209]=30'd475492838;
array[17210]=30'd461875644;
array[17211]=30'd414702010;
array[17212]=30'd359126474;
array[17213]=30'd422024669;
array[17214]=30'd597116464;
array[17215]=30'd883367490;
array[17216]=30'd855016073;
array[17217]=30'd695644807;
array[17218]=30'd695644807;
array[17219]=30'd855016073;
array[17220]=30'd855016073;
array[17221]=30'd855016073;
array[17222]=30'd855016073;
array[17223]=30'd855016073;
array[17224]=30'd583395966;
array[17225]=30'd637892242;
array[17226]=30'd601183923;
array[17227]=30'd463850128;
array[17228]=30'd637892242;
array[17229]=30'd568787568;
array[17230]=30'd842497613;
array[17231]=30'd804744750;
array[17232]=30'd504834577;
array[17233]=30'd396849695;
array[17234]=30'd722945572;
array[17235]=30'd768057919;
array[17236]=30'd555187752;
array[17237]=30'd468145703;
array[17238]=30'd959930934;
array[17239]=30'd979844654;
array[17240]=30'd979844654;
array[17241]=30'd959930934;
array[17242]=30'd959930934;
array[17243]=30'd959930934;
array[17244]=30'd959930934;
array[17245]=30'd650619404;
array[17246]=30'd333946399;
array[17247]=30'd597116464;
array[17248]=30'd679961142;
array[17249]=30'd468145703;
array[17250]=30'd258428439;
array[17251]=30'd504834577;
array[17252]=30'd679961142;
array[17253]=30'd893852174;
array[17254]=30'd959930934;
array[17255]=30'd916919852;
array[17256]=30'd792119862;
array[17257]=30'd583395966;
array[17258]=30'd637892242;
array[17259]=30'd452327079;
array[17260]=30'd646252225;
array[17261]=30'd646252225;
array[17262]=30'd601183923;
array[17263]=30'd556097214;
array[17264]=30'd646252225;
array[17265]=30'd548775573;
array[17266]=30'd879170165;
array[17267]=30'd879170165;
array[17268]=30'd879170165;
array[17269]=30'd879170165;
array[17270]=30'd879170165;
array[17271]=30'd879170165;
array[17272]=30'd900141674;
array[17273]=30'd900141674;
array[17274]=30'd879170165;
array[17275]=30'd879170165;
array[17276]=30'd879170165;
array[17277]=30'd879170165;
array[17278]=30'd855016073;
array[17279]=30'd855016073;
array[17280]=30'd855016073;
array[17281]=30'd855016073;
array[17282]=30'd855016073;
array[17283]=30'd879170165;
array[17284]=30'd879170165;
array[17285]=30'd879170165;
array[17286]=30'd879170165;
array[17287]=30'd879170165;
array[17288]=30'd879170165;
array[17289]=30'd922198619;
array[17290]=30'd996656669;
array[17291]=30'd894969309;
array[17292]=30'd785935846;
array[17293]=30'd855121400;
array[17294]=30'd983041534;
array[17295]=30'd872938009;
array[17296]=30'd414702010;
array[17297]=30'd479712691;
array[17298]=30'd490193319;
array[17299]=30'd490193319;
array[17300]=30'd479712691;
array[17301]=30'd461875644;
array[17302]=30'd525848010;
array[17303]=30'd422024669;
array[17304]=30'd461875644;
array[17305]=30'd461875644;
array[17306]=30'd448250284;
array[17307]=30'd359126474;
array[17308]=30'd359126474;
array[17309]=30'd341278169;
array[17310]=30'd722945572;
array[17311]=30'd883367490;
array[17312]=30'd855016073;
array[17313]=30'd855016073;
array[17314]=30'd779516542;
array[17315]=30'd695644807;
array[17316]=30'd816210575;
array[17317]=30'd855016073;
array[17318]=30'd855016073;
array[17319]=30'd855016073;
array[17320]=30'd624350812;
array[17321]=30'd614845038;
array[17322]=30'd559303301;
array[17323]=30'd337060463;
array[17324]=30'd417795660;
array[17325]=30'd417795660;
array[17326]=30'd804744750;
array[17327]=30'd352806463;
array[17328]=30'd613923367;
array[17329]=30'd916919852;
array[17330]=30'd959930934;
array[17331]=30'd959930934;
array[17332]=30'd959930934;
array[17333]=30'd883367490;
array[17334]=30'd959930934;
array[17335]=30'd959930934;
array[17336]=30'd979844654;
array[17337]=30'd959930934;
array[17338]=30'd959930934;
array[17339]=30'd959930934;
array[17340]=30'd959930934;
array[17341]=30'd859252262;
array[17342]=30'd916919852;
array[17343]=30'd959930934;
array[17344]=30'd959930934;
array[17345]=30'd959930934;
array[17346]=30'd804744750;
array[17347]=30'd468145703;
array[17348]=30'd294108730;
array[17349]=30'd804744750;
array[17350]=30'd959930934;
array[17351]=30'd941029952;
array[17352]=30'd751243845;
array[17353]=30'd614845038;
array[17354]=30'd637892242;
array[17355]=30'd427157133;
array[17356]=30'd518350503;
array[17357]=30'd646252225;
array[17358]=30'd556097214;
array[17359]=30'd601183923;
array[17360]=30'd668323493;
array[17361]=30'd624350812;
array[17362]=30'd941029952;
array[17363]=30'd883367490;
array[17364]=30'd883367490;
array[17365]=30'd916919852;
array[17366]=30'd936883742;
array[17367]=30'd936883742;
array[17368]=30'd960978443;
array[17369]=30'd960978443;
array[17370]=30'd979844654;
array[17371]=30'd941029952;
array[17372]=30'd879170165;
array[17373]=30'd879170165;
array[17374]=30'd879170165;
array[17375]=30'd855016073;
array[17376]=30'd855016073;
array[17377]=30'd855016073;
array[17378]=30'd855016073;
array[17379]=30'd879170165;
array[17380]=30'd879170165;
array[17381]=30'd879170165;
array[17382]=30'd879170165;
array[17383]=30'd879170165;
array[17384]=30'd900141674;
array[17385]=30'd959930934;
array[17386]=30'd898098744;
array[17387]=30'd777516526;
array[17388]=30'd815247846;
array[17389]=30'd893852174;
array[17390]=30'd996656669;
array[17391]=30'd855121400;
array[17392]=30'd414702010;
array[17393]=30'd490193319;
array[17394]=30'd490193319;
array[17395]=30'd479712691;
array[17396]=30'd448250284;
array[17397]=30'd394764738;
array[17398]=30'd414702010;
array[17399]=30'd461875644;
array[17400]=30'd479712691;
array[17401]=30'd479712691;
array[17402]=30'd448250284;
array[17403]=30'd448250284;
array[17404]=30'd475492838;
array[17405]=30'd722945572;
array[17406]=30'd665233987;
array[17407]=30'd794239590;
array[17408]=30'd855016073;
array[17409]=30'd855016073;
array[17410]=30'd855016073;
array[17411]=30'd855016073;
array[17412]=30'd730239616;
array[17413]=30'd779516542;
array[17414]=30'd879170165;
array[17415]=30'd879170165;
array[17416]=30'd624350812;
array[17417]=30'd417795660;
array[17418]=30'd396849695;
array[17419]=30'd475492838;
array[17420]=30'd475492838;
array[17421]=30'd442989058;
array[17422]=30'd300376570;
array[17423]=30'd617028085;
array[17424]=30'd959930934;
array[17425]=30'd979844654;
array[17426]=30'd959930934;
array[17427]=30'd959930934;
array[17428]=30'd959930934;
array[17429]=30'd959930934;
array[17430]=30'd959930934;
array[17431]=30'd959930934;
array[17432]=30'd959930934;
array[17433]=30'd959930934;
array[17434]=30'd979844654;
array[17435]=30'd959930934;
array[17436]=30'd959930934;
array[17437]=30'd979844654;
array[17438]=30'd959930934;
array[17439]=30'd959930934;
array[17440]=30'd959930934;
array[17441]=30'd959930934;
array[17442]=30'd959930934;
array[17443]=30'd916919852;
array[17444]=30'd555187752;
array[17445]=30'd396849695;
array[17446]=30'd959930934;
array[17447]=30'd941029952;
array[17448]=30'd665233987;
array[17449]=30'd614845038;
array[17450]=30'd601183923;
array[17451]=30'd394645149;
array[17452]=30'd556097214;
array[17453]=30'd646252225;
array[17454]=30'd518350503;
array[17455]=30'd601183923;
array[17456]=30'd611709603;
array[17457]=30'd671568495;
array[17458]=30'd936883742;
array[17459]=30'd872938009;
array[17460]=30'd855121400;
array[17461]=30'd832062938;
array[17462]=30'd785935846;
array[17463]=30'd767069629;
array[17464]=30'd809003452;
array[17465]=30'd809003452;
array[17466]=30'd928507337;
array[17467]=30'd960978443;
array[17468]=30'd916919852;
array[17469]=30'd879170165;
array[17470]=30'd879170165;
array[17471]=30'd855016073;
array[17472]=30'd855016073;
array[17473]=30'd879170165;
array[17474]=30'd879170165;
array[17475]=30'd879170165;
array[17476]=30'd879170165;
array[17477]=30'd879170165;
array[17478]=30'd879170165;
array[17479]=30'd879170165;
array[17480]=30'd879170165;
array[17481]=30'd922198619;
array[17482]=30'd842497613;
array[17483]=30'd839346691;
array[17484]=30'd893852174;
array[17485]=30'd916919852;
array[17486]=30'd959930934;
array[17487]=30'd832062938;
array[17488]=30'd461875644;
array[17489]=30'd479712691;
array[17490]=30'd490193319;
array[17491]=30'd479712691;
array[17492]=30'd414702010;
array[17493]=30'd414702010;
array[17494]=30'd479712691;
array[17495]=30'd479712691;
array[17496]=30'd479712691;
array[17497]=30'd479712691;
array[17498]=30'd448250284;
array[17499]=30'd475492838;
array[17500]=30'd792119862;
array[17501]=30'd883367490;
array[17502]=30'd824630873;
array[17503]=30'd730239616;
array[17504]=30'd779516542;
array[17505]=30'd879170165;
array[17506]=30'd879170165;
array[17507]=30'd879170165;
array[17508]=30'd879170165;
array[17509]=30'd794239590;
array[17510]=30'd671568495;
array[17511]=30'd751243845;
array[17512]=30'd468145703;
array[17513]=30'd442989058;
array[17514]=30'd461875644;
array[17515]=30'd461875644;
array[17516]=30'd448250284;
array[17517]=30'd372750770;
array[17518]=30'd554095113;
array[17519]=30'd761730564;
array[17520]=30'd959930934;
array[17521]=30'd959930934;
array[17522]=30'd959930934;
array[17523]=30'd959930934;
array[17524]=30'd959930934;
array[17525]=30'd959930934;
array[17526]=30'd959930934;
array[17527]=30'd959930934;
array[17528]=30'd959930934;
array[17529]=30'd959930934;
array[17530]=30'd959930934;
array[17531]=30'd959930934;
array[17532]=30'd959930934;
array[17533]=30'd959930934;
array[17534]=30'd959930934;
array[17535]=30'd959930934;
array[17536]=30'd959930934;
array[17537]=30'd959930934;
array[17538]=30'd959930934;
array[17539]=30'd959930934;
array[17540]=30'd941029952;
array[17541]=30'd804744750;
array[17542]=30'd959930934;
array[17543]=30'd941029952;
array[17544]=30'd624350812;
array[17545]=30'd637892242;
array[17546]=30'd601183923;
array[17547]=30'd394645149;
array[17548]=30'd601183923;
array[17549]=30'd646252225;
array[17550]=30'd486895284;
array[17551]=30'd668323493;
array[17552]=30'd556097214;
array[17553]=30'd751243845;
array[17554]=30'd820526616;
array[17555]=30'd785935846;
array[17556]=30'd767069629;
array[17557]=30'd767069629;
array[17558]=30'd809003452;
array[17559]=30'd809003452;
array[17560]=30'd849905057;
array[17561]=30'd829990281;
array[17562]=30'd792242589;
array[17563]=30'd928507337;
array[17564]=30'd960978443;
array[17565]=30'd883367490;
array[17566]=30'd879170165;
array[17567]=30'd855016073;
array[17568]=30'd879170165;
array[17569]=30'd879170165;
array[17570]=30'd879170165;
array[17571]=30'd879170165;
array[17572]=30'd879170165;
array[17573]=30'd879170165;
array[17574]=30'd879170165;
array[17575]=30'd879170165;
array[17576]=30'd879170165;
array[17577]=30'd900141674;
array[17578]=30'd883367490;
array[17579]=30'd883367490;
array[17580]=30'd879170165;
array[17581]=30'd900141674;
array[17582]=30'd898098744;
array[17583]=30'd777516526;
array[17584]=30'd441989592;
array[17585]=30'd490193319;
array[17586]=30'd490193319;
array[17587]=30'd479712691;
array[17588]=30'd372750770;
array[17589]=30'd479712691;
array[17590]=30'd479712691;
array[17591]=30'd479712691;
array[17592]=30'd479712691;
array[17593]=30'd461875644;
array[17594]=30'd525848010;
array[17595]=30'd804744750;
array[17596]=30'd883367490;
array[17597]=30'd879170165;
array[17598]=30'd879170165;
array[17599]=30'd879170165;
array[17600]=30'd779516542;
array[17601]=30'd730239616;
array[17602]=30'd879170165;
array[17603]=30'd879170165;
array[17604]=30'd879170165;
array[17605]=30'd824630873;
array[17606]=30'd527922743;
array[17607]=30'd333946399;
array[17608]=30'd475492838;
array[17609]=30'd479712691;
array[17610]=30'd448250284;
array[17611]=30'd394764738;
array[17612]=30'd372750770;
array[17613]=30'd359126474;
array[17614]=30'd684132856;
array[17615]=30'd804744750;
array[17616]=30'd679961142;
array[17617]=30'd916919852;
array[17618]=30'd941029952;
array[17619]=30'd916919852;
array[17620]=30'd959930934;
array[17621]=30'd959930934;
array[17622]=30'd959930934;
array[17623]=30'd959930934;
array[17624]=30'd959930934;
array[17625]=30'd959930934;
array[17626]=30'd959930934;
array[17627]=30'd959930934;
array[17628]=30'd959930934;
array[17629]=30'd959930934;
array[17630]=30'd959930934;
array[17631]=30'd959930934;
array[17632]=30'd941029952;
array[17633]=30'd883367490;
array[17634]=30'd959930934;
array[17635]=30'd941029952;
array[17636]=30'd883367490;
array[17637]=30'd959930934;
array[17638]=30'd941029952;
array[17639]=30'd916919852;
array[17640]=30'd527849061;
array[17641]=30'd637892242;
array[17642]=30'd556097214;
array[17643]=30'd394645149;
array[17644]=30'd601183923;
array[17645]=30'd646252225;
array[17646]=30'd518350503;
array[17647]=30'd646252225;
array[17648]=30'd548775573;
array[17649]=30'd802671197;
array[17650]=30'd820526616;
array[17651]=30'd785935846;
array[17652]=30'd832062938;
array[17653]=30'd894969309;
array[17654]=30'd928507337;
array[17655]=30'd893925805;
array[17656]=30'd849905057;
array[17657]=30'd876132737;
array[17658]=30'd829990281;
array[17659]=30'd809003452;
array[17660]=30'd948416998;
array[17661]=30'd916919852;
array[17662]=30'd883367490;
array[17663]=30'd855016073;
array[17664]=30'd879170165;
array[17665]=30'd879170165;
array[17666]=30'd879170165;
array[17667]=30'd879170165;
array[17668]=30'd879170165;
array[17669]=30'd879170165;
array[17670]=30'd879170165;
array[17671]=30'd879170165;
array[17672]=30'd879170165;
array[17673]=30'd879170165;
array[17674]=30'd879170165;
array[17675]=30'd879170165;
array[17676]=30'd879170165;
array[17677]=30'd879170165;
array[17678]=30'd900141674;
array[17679]=30'd820526616;
array[17680]=30'd461903352;
array[17681]=30'd479712691;
array[17682]=30'd479712691;
array[17683]=30'd479712691;
array[17684]=30'd448250284;
array[17685]=30'd490193319;
array[17686]=30'd479712691;
array[17687]=30'd461875644;
array[17688]=30'd448250284;
array[17689]=30'd571957759;
array[17690]=30'd859252262;
array[17691]=30'd883367490;
array[17692]=30'd879170165;
array[17693]=30'd879170165;
array[17694]=30'd879170165;
array[17695]=30'd879170165;
array[17696]=30'd879170165;
array[17697]=30'd816210575;
array[17698]=30'd730239616;
array[17699]=30'd879170165;
array[17700]=30'd824630873;
array[17701]=30'd597116464;
array[17702]=30'd442989058;
array[17703]=30'd475492838;
array[17704]=30'd394764738;
array[17705]=30'd394764738;
array[17706]=30'd394764738;
array[17707]=30'd414702010;
array[17708]=30'd372750770;
array[17709]=30'd341278169;
array[17710]=30'd839346691;
array[17711]=30'd959930934;
array[17712]=30'd768057919;
array[17713]=30'd804744750;
array[17714]=30'd959930934;
array[17715]=30'd959930934;
array[17716]=30'd959930934;
array[17717]=30'd959930934;
array[17718]=30'd959930934;
array[17719]=30'd959930934;
array[17720]=30'd959930934;
array[17721]=30'd959930934;
array[17722]=30'd959930934;
array[17723]=30'd959930934;
array[17724]=30'd959930934;
array[17725]=30'd959930934;
array[17726]=30'd959930934;
array[17727]=30'd959930934;
array[17728]=30'd916919852;
array[17729]=30'd941029952;
array[17730]=30'd959930934;
array[17731]=30'd883367490;
array[17732]=30'd941029952;
array[17733]=30'd959930934;
array[17734]=30'd842497613;
array[17735]=30'd859252262;
array[17736]=30'd527849061;
array[17737]=30'd637892242;
array[17738]=30'd518350503;
array[17739]=30'd497425057;
array[17740]=30'd668323493;
array[17741]=30'd556097214;
array[17742]=30'd556097214;
array[17743]=30'd646252225;
array[17744]=30'd559303301;
array[17745]=30'd857217603;
array[17746]=30'd785935846;
array[17747]=30'd832062938;
array[17748]=30'd894969309;
array[17749]=30'd832062938;
array[17750]=30'd785935846;
array[17751]=30'd767069629;
array[17752]=30'd778590630;
array[17753]=30'd766030218;
array[17754]=30'd829990281;
array[17755]=30'd792242589;
array[17756]=30'd893925805;
array[17757]=30'd960978443;
array[17758]=30'd883367490;
array[17759]=30'd855016073;
array[17760]=30'd900141674;
array[17761]=30'd883367490;
array[17762]=30'd883367490;
array[17763]=30'd883367490;
array[17764]=30'd900141674;
array[17765]=30'd879170165;
array[17766]=30'd879170165;
array[17767]=30'd879170165;
array[17768]=30'd879170165;
array[17769]=30'd879170165;
array[17770]=30'd879170165;
array[17771]=30'd900141674;
array[17772]=30'd879170165;
array[17773]=30'd879170165;
array[17774]=30'd879170165;
array[17775]=30'd857217603;
array[17776]=30'd483930653;
array[17777]=30'd492300766;
array[17778]=30'd490193319;
array[17779]=30'd479712691;
array[17780]=30'd479712691;
array[17781]=30'd479712691;
array[17782]=30'd461875644;
array[17783]=30'd422024669;
array[17784]=30'd650619404;
array[17785]=30'd859252262;
array[17786]=30'd879170165;
array[17787]=30'd879170165;
array[17788]=30'd879170165;
array[17789]=30'd879170165;
array[17790]=30'd879170165;
array[17791]=30'd879170165;
array[17792]=30'd879170165;
array[17793]=30'd879170165;
array[17794]=30'd824630873;
array[17795]=30'd597116464;
array[17796]=30'd504834577;
array[17797]=30'd475492838;
array[17798]=30'd479712691;
array[17799]=30'd461875644;
array[17800]=30'd448250284;
array[17801]=30'd359126474;
array[17802]=30'd448250284;
array[17803]=30'd448250284;
array[17804]=30'd414702010;
array[17805]=30'd422024669;
array[17806]=30'd804744750;
array[17807]=30'd959930934;
array[17808]=30'd959930934;
array[17809]=30'd768057919;
array[17810]=30'd916919852;
array[17811]=30'd959930934;
array[17812]=30'd959930934;
array[17813]=30'd959930934;
array[17814]=30'd959930934;
array[17815]=30'd959930934;
array[17816]=30'd959930934;
array[17817]=30'd979844654;
array[17818]=30'd979844654;
array[17819]=30'd959930934;
array[17820]=30'd959930934;
array[17821]=30'd959930934;
array[17822]=30'd959930934;
array[17823]=30'd959930934;
array[17824]=30'd941029952;
array[17825]=30'd959930934;
array[17826]=30'd959930934;
array[17827]=30'd959930934;
array[17828]=30'd959930934;
array[17829]=30'd941029952;
array[17830]=30'd941029952;
array[17831]=30'd792119862;
array[17832]=30'd559303301;
array[17833]=30'd637892242;
array[17834]=30'd463850128;
array[17835]=30'd556097214;
array[17836]=30'd668323493;
array[17837]=30'd518350503;
array[17838]=30'd611709603;
array[17839]=30'd601183923;
array[17840]=30'd651585154;
array[17841]=30'd820526616;
array[17842]=30'd785935846;
array[17843]=30'd894969309;
array[17844]=30'd872938009;
array[17845]=30'd785935846;
array[17846]=30'd809003452;
array[17847]=30'd893925805;
array[17848]=30'd849905057;
array[17849]=30'd778590630;
array[17850]=30'd849905057;
array[17851]=30'd876132737;
array[17852]=30'd809003452;
array[17853]=30'd948416998;
array[17854]=30'd883367490;
array[17855]=30'd879170165;
array[17856]=30'd900141674;
array[17857]=30'd893852174;
array[17858]=30'd871846383;
array[17859]=30'd893852174;
array[17860]=30'd883367490;
array[17861]=30'd883367490;
array[17862]=30'd879170165;
array[17863]=30'd879170165;
array[17864]=30'd879170165;
array[17865]=30'd879170165;
array[17866]=30'd900141674;
array[17867]=30'd900141674;
array[17868]=30'd879170165;
array[17869]=30'd879170165;
array[17870]=30'd879170165;
array[17871]=30'd879170165;
array[17872]=30'd468145703;
array[17873]=30'd492300766;
array[17874]=30'd479712691;
array[17875]=30'd479712691;
array[17876]=30'd479712691;
array[17877]=30'd448250284;
array[17878]=30'd479712691;
array[17879]=30'd761730564;
array[17880]=30'd859252262;
array[17881]=30'd879170165;
array[17882]=30'd879170165;
array[17883]=30'd879170165;
array[17884]=30'd879170165;
array[17885]=30'd879170165;
array[17886]=30'd879170165;
array[17887]=30'd879170165;
array[17888]=30'd879170165;
array[17889]=30'd879170165;
array[17890]=30'd794239590;
array[17891]=30'd468145703;
array[17892]=30'd387463674;
array[17893]=30'd461875644;
array[17894]=30'd479712691;
array[17895]=30'd479712691;
array[17896]=30'd479712691;
array[17897]=30'd414702010;
array[17898]=30'd394764738;
array[17899]=30'd479712691;
array[17900]=30'd414702010;
array[17901]=30'd504834577;
array[17902]=30'd893852174;
array[17903]=30'd959930934;
array[17904]=30'd959930934;
array[17905]=30'd941029952;
array[17906]=30'd722945572;
array[17907]=30'd597116464;
array[17908]=30'd597116464;
array[17909]=30'd641176139;
array[17910]=30'd679961142;
array[17911]=30'd751243845;
array[17912]=30'd804744750;
array[17913]=30'd804744750;
array[17914]=30'd804744750;
array[17915]=30'd804744750;
array[17916]=30'd751243845;
array[17917]=30'd722945572;
array[17918]=30'd679961142;
array[17919]=30'd597116464;
array[17920]=30'd527922743;
array[17921]=30'd679961142;
array[17922]=30'd959930934;
array[17923]=30'd959930934;
array[17924]=30'd959930934;
array[17925]=30'd959930934;
array[17926]=30'd941029952;
array[17927]=30'd751243845;
array[17928]=30'd614845038;
array[17929]=30'd601183923;
array[17930]=30'd427157133;
array[17931]=30'd601183923;
array[17932]=30'd601183923;
array[17933]=30'd463850128;
array[17934]=30'd637892242;
array[17935]=30'd583395966;
array[17936]=30'd707208791;
array[17937]=30'd820526616;
array[17938]=30'd785935846;
array[17939]=30'd894969309;
array[17940]=30'd872938009;
array[17941]=30'd785935846;
array[17942]=30'd809003452;
array[17943]=30'd977825191;
array[17944]=30'd893925805;
array[17945]=30'd809003452;
array[17946]=30'd792242589;
array[17947]=30'd908629408;
array[17948]=30'd778590630;
array[17949]=30'd894969309;
array[17950]=30'd916919852;
array[17951]=30'd879170165;
array[17952]=30'd857217603;
array[17953]=30'd855121400;
array[17954]=30'd871846383;
array[17955]=30'd871846383;
array[17956]=30'd893852174;
array[17957]=30'd883367490;
array[17958]=30'd900141674;
array[17959]=30'd900141674;
array[17960]=30'd900141674;
array[17961]=30'd879170165;
array[17962]=30'd879170165;
array[17963]=30'd900141674;
array[17964]=30'd879170165;
array[17965]=30'd879170165;
array[17966]=30'd879170165;
array[17967]=30'd879170165;
array[17968]=30'd527922743;
array[17969]=30'd492300766;
array[17970]=30'd479712691;
array[17971]=30'd461875644;
array[17972]=30'd422024669;
array[17973]=30'd617028085;
array[17974]=30'd804744750;
array[17975]=30'd883367490;
array[17976]=30'd879170165;
array[17977]=30'd879170165;
array[17978]=30'd879170165;
array[17979]=30'd879170165;
array[17980]=30'd879170165;
array[17981]=30'd879170165;
array[17982]=30'd879170165;
array[17983]=30'd879170165;
array[17984]=30'd879170165;
array[17985]=30'd824630873;
array[17986]=30'd527922743;
array[17987]=30'd461903352;
array[17988]=30'd461875644;
array[17989]=30'd414702010;
array[17990]=30'd479712691;
array[17991]=30'd479712691;
array[17992]=30'd479712691;
array[17993]=30'd461875644;
array[17994]=30'd359126474;
array[17995]=30'd341278169;
array[17996]=30'd442989058;
array[17997]=30'd804744750;
array[17998]=30'd959930934;
array[17999]=30'd959930934;
array[18000]=30'd959930934;
array[18001]=30'd959930934;
array[18002]=30'd883367490;
array[18003]=30'd417795660;
array[18004]=30'd352806463;
array[18005]=30'd385301087;
array[18006]=30'd385301087;
array[18007]=30'd385301087;
array[18008]=30'd385301087;
array[18009]=30'd385301087;
array[18010]=30'd385301087;
array[18011]=30'd385301087;
array[18012]=30'd385301087;
array[18013]=30'd385301087;
array[18014]=30'd385301087;
array[18015]=30'd385301087;
array[18016]=30'd385301087;
array[18017]=30'd468145703;
array[18018]=30'd959930934;
array[18019]=30'd959930934;
array[18020]=30'd959930934;
array[18021]=30'd959930934;
array[18022]=30'd941029952;
array[18023]=30'd624350812;
array[18024]=30'd637892242;
array[18025]=30'd637892242;
array[18026]=30'd497425057;
array[18027]=30'd637892242;
array[18028]=30'd556097214;
array[18029]=30'd463850128;
array[18030]=30'd668323493;
array[18031]=30'd548775573;
array[18032]=30'd794239590;
array[18033]=30'd820526616;
array[18034]=30'd767069629;
array[18035]=30'd928507337;
array[18036]=30'd893852174;
array[18037]=30'd820526616;
array[18038]=30'd767069629;
array[18039]=30'd945318330;
array[18040]=30'd871910847;
array[18041]=30'd809003452;
array[18042]=30'd792242589;
array[18043]=30'd908629408;
array[18044]=30'd778590630;
array[18045]=30'd871910847;
array[18046]=30'd893852174;
array[18047]=30'd879170165;
array[18048]=30'd872938009;
array[18049]=30'd855121400;
array[18050]=30'd855121400;
array[18051]=30'd871846383;
array[18052]=30'd859252262;
array[18053]=30'd883367490;
array[18054]=30'd900141674;
array[18055]=30'd900141674;
array[18056]=30'd900141674;
array[18057]=30'd900141674;
array[18058]=30'd879170165;
array[18059]=30'd879170165;
array[18060]=30'd879170165;
array[18061]=30'd900141674;
array[18062]=30'd879170165;
array[18063]=30'd879170165;
array[18064]=30'd571952708;
array[18065]=30'd492300766;
array[18066]=30'd479712691;
array[18067]=30'd414702010;
array[18068]=30'd694663659;
array[18069]=30'd883367490;
array[18070]=30'd883367490;
array[18071]=30'd900141674;
array[18072]=30'd900141674;
array[18073]=30'd879170165;
array[18074]=30'd879170165;
array[18075]=30'd900141674;
array[18076]=30'd879170165;
array[18077]=30'd879170165;
array[18078]=30'd879170165;
array[18079]=30'd879170165;
array[18080]=30'd842497613;
array[18081]=30'd555187752;
array[18082]=30'd492300766;
array[18083]=30'd492300766;
array[18084]=30'd479712691;
array[18085]=30'd448250284;
array[18086]=30'd394764738;
array[18087]=30'd461875644;
array[18088]=30'd414702010;
array[18089]=30'd422024669;
array[18090]=30'd396849695;
array[18091]=30'd378982955;
array[18092]=30'd583428668;
array[18093]=30'd665233987;
array[18094]=30'd941029952;
array[18095]=30'd959930934;
array[18096]=30'd959930934;
array[18097]=30'd959930934;
array[18098]=30'd959930934;
array[18099]=30'd722945572;
array[18100]=30'd352806463;
array[18101]=30'd385301087;
array[18102]=30'd385301087;
array[18103]=30'd385301087;
array[18104]=30'd385301087;
array[18105]=30'd385301087;
array[18106]=30'd385301087;
array[18107]=30'd385301087;
array[18108]=30'd385301087;
array[18109]=30'd385301087;
array[18110]=30'd385301087;
array[18111]=30'd385301087;
array[18112]=30'd385301087;
array[18113]=30'd597116464;
array[18114]=30'd959930934;
array[18115]=30'd959930934;
array[18116]=30'd941029952;
array[18117]=30'd941029952;
array[18118]=30'd916919852;
array[18119]=30'd557205073;
array[18120]=30'd637892242;
array[18121]=30'd548775573;
array[18122]=30'd601183923;
array[18123]=30'd601183923;
array[18124]=30'd463850128;
array[18125]=30'd523632283;
array[18126]=30'd668323493;
array[18127]=30'd559303301;
array[18128]=30'd883367490;
array[18129]=30'd820526616;
array[18130]=30'd809003452;
array[18131]=30'd948416998;
array[18132]=30'd872938009;
array[18133]=30'd820526616;
array[18134]=30'd785935846;
array[18135]=30'd893925805;
array[18136]=30'd871910847;
array[18137]=30'd767069629;
array[18138]=30'd792242589;
array[18139]=30'd829990281;
array[18140]=30'd778590630;
array[18141]=30'd894969309;
array[18142]=30'd859252262;
array[18143]=30'd879170165;
array[18144]=30'd872938009;
array[18145]=30'd855121400;
array[18146]=30'd894969309;
array[18147]=30'd871846383;
array[18148]=30'd893852174;
array[18149]=30'd900141674;
array[18150]=30'd900141674;
array[18151]=30'd900141674;
array[18152]=30'd900141674;
array[18153]=30'd900141674;
array[18154]=30'd900141674;
array[18155]=30'd900141674;
array[18156]=30'd900141674;
array[18157]=30'd900141674;
array[18158]=30'd879170165;
array[18159]=30'd900141674;
array[18160]=30'd641176139;
array[18161]=30'd461903352;
array[18162]=30'd479712691;
array[18163]=30'd525848010;
array[18164]=30'd859252262;
array[18165]=30'd883367490;
array[18166]=30'd900141674;
array[18167]=30'd900141674;
array[18168]=30'd900141674;
array[18169]=30'd900141674;
array[18170]=30'd900141674;
array[18171]=30'd900141674;
array[18172]=30'd879170165;
array[18173]=30'd879170165;
array[18174]=30'd879170165;
array[18175]=30'd879170165;
array[18176]=30'd597116464;
array[18177]=30'd461903352;
array[18178]=30'd479712691;
array[18179]=30'd479712691;
array[18180]=30'd479712691;
array[18181]=30'd479712691;
array[18182]=30'd359126474;
array[18183]=30'd394764738;
array[18184]=30'd684132856;
array[18185]=30'd792119862;
array[18186]=30'd484882002;
array[18187]=30'd406210138;
array[18188]=30'd484816502;
array[18189]=30'd559303301;
array[18190]=30'd824630873;
array[18191]=30'd941029952;
array[18192]=30'd959930934;
array[18193]=30'd959930934;
array[18194]=30'd959930934;
array[18195]=30'd916919852;
array[18196]=30'd468145703;
array[18197]=30'd385301087;
array[18198]=30'd417795660;
array[18199]=30'd457612903;
array[18200]=30'd484882002;
array[18201]=30'd457612903;
array[18202]=30'd457612903;
array[18203]=30'd457612903;
array[18204]=30'd417795660;
array[18205]=30'd385301087;
array[18206]=30'd385301087;
array[18207]=30'd385301087;
array[18208]=30'd417795660;
array[18209]=30'd859252262;
array[18210]=30'd959930934;
array[18211]=30'd959930934;
array[18212]=30'd959930934;
array[18213]=30'd941029952;
array[18214]=30'd883367490;
array[18215]=30'd527849061;
array[18216]=30'd637892242;
array[18217]=30'd444947126;
array[18218]=30'd668323493;
array[18219]=30'd556097214;
array[18220]=30'd324381369;
array[18221]=30'd611709603;
array[18222]=30'd637892242;
array[18223]=30'd593953387;
array[18224]=30'd900141674;
array[18225]=30'd820526616;
array[18226]=30'd785935846;
array[18227]=30'd965227994;
array[18228]=30'd936883742;
array[18229]=30'd820526616;
array[18230]=30'd785935846;
array[18231]=30'd871910847;
array[18232]=30'd977825191;
array[18233]=30'd945318330;
array[18234]=30'd908629408;
array[18235]=30'd809003452;
array[18236]=30'd809003452;
array[18237]=30'd916977147;
array[18238]=30'd883367490;
array[18239]=30'd879170165;
array[18240]=30'd872938009;
array[18241]=30'd872938009;
array[18242]=30'd893852174;
array[18243]=30'd893852174;
array[18244]=30'd883367490;
array[18245]=30'd900141674;
array[18246]=30'd900141674;
array[18247]=30'd900141674;
array[18248]=30'd900141674;
array[18249]=30'd900141674;
array[18250]=30'd900141674;
array[18251]=30'd900141674;
array[18252]=30'd900141674;
array[18253]=30'd900141674;
array[18254]=30'd879170165;
array[18255]=30'd900141674;
array[18256]=30'd679961142;
array[18257]=30'd475492838;
array[18258]=30'd479712691;
array[18259]=30'd475492838;
array[18260]=30'd883367490;
array[18261]=30'd900141674;
array[18262]=30'd900141674;
array[18263]=30'd900141674;
array[18264]=30'd900141674;
array[18265]=30'd900141674;
array[18266]=30'd900141674;
array[18267]=30'd900141674;
array[18268]=30'd900141674;
array[18269]=30'd900141674;
array[18270]=30'd900141674;
array[18271]=30'd679961142;
array[18272]=30'd442989058;
array[18273]=30'd479712691;
array[18274]=30'd490193319;
array[18275]=30'd479712691;
array[18276]=30'd461875644;
array[18277]=30'd461875644;
array[18278]=30'd619182551;
array[18279]=30'd617028085;
array[18280]=30'd804744750;
array[18281]=30'd883367490;
array[18282]=30'd484882002;
array[18283]=30'd406210138;
array[18284]=30'd527849061;
array[18285]=30'd484816502;
array[18286]=30'd457612903;
array[18287]=30'd751243845;
array[18288]=30'd941029952;
array[18289]=30'd959930934;
array[18290]=30'd959930934;
array[18291]=30'd959930934;
array[18292]=30'd859252262;
array[18293]=30'd417795660;
array[18294]=30'd593953387;
array[18295]=30'd624350812;
array[18296]=30'd624350812;
array[18297]=30'd624350812;
array[18298]=30'd624350812;
array[18299]=30'd593953387;
array[18300]=30'd593953387;
array[18301]=30'd548890196;
array[18302]=30'd484882002;
array[18303]=30'd417795660;
array[18304]=30'd804744750;
array[18305]=30'd959930934;
array[18306]=30'd959930934;
array[18307]=30'd959930934;
array[18308]=30'd941029952;
array[18309]=30'd941029952;
array[18310]=30'd624350812;
array[18311]=30'd583395966;
array[18312]=30'd548775573;
array[18313]=30'd556097214;
array[18314]=30'd601183923;
array[18315]=30'd452327079;
array[18316]=30'd394645149;
array[18317]=30'd611709603;
array[18318]=30'd611709603;
array[18319]=30'd695644807;
array[18320]=30'd900141674;
array[18321]=30'd857217603;
array[18322]=30'd785935846;
array[18323]=30'd928507337;
array[18324]=30'd983041534;
array[18325]=30'd916977147;
array[18326]=30'd785935846;
array[18327]=30'd767069629;
array[18328]=30'd871910847;
array[18329]=30'd945318330;
array[18330]=30'd893925805;
array[18331]=30'd778590630;
array[18332]=30'd815247846;
array[18333]=30'd893852174;
array[18334]=30'd883367490;
array[18335]=30'd879170165;
array[18336]=30'd900141674;
array[18337]=30'd898098744;
array[18338]=30'd883367490;
array[18339]=30'd883367490;
array[18340]=30'd900141674;
array[18341]=30'd900141674;
array[18342]=30'd900141674;
array[18343]=30'd900141674;
array[18344]=30'd900141674;
array[18345]=30'd900141674;
array[18346]=30'd900141674;
array[18347]=30'd900141674;
array[18348]=30'd900141674;
array[18349]=30'd879170165;
array[18350]=30'd900141674;
array[18351]=30'd879170165;
array[18352]=30'd751243845;
array[18353]=30'd442989058;
array[18354]=30'd479712691;
array[18355]=30'd442989058;
array[18356]=30'd859252262;
array[18357]=30'd900141674;
array[18358]=30'd900141674;
array[18359]=30'd900141674;
array[18360]=30'd900141674;
array[18361]=30'd900141674;
array[18362]=30'd900141674;
array[18363]=30'd900141674;
array[18364]=30'd900141674;
array[18365]=30'd900141674;
array[18366]=30'd751243845;
array[18367]=30'd468145703;
array[18368]=30'd492300766;
array[18369]=30'd490193319;
array[18370]=30'd479712691;
array[18371]=30'd414702010;
array[18372]=30'd414702010;
array[18373]=30'd619182551;
array[18374]=30'd777516526;
array[18375]=30'd597116464;
array[18376]=30'd527922743;
array[18377]=30'd679961142;
array[18378]=30'd449215039;
array[18379]=30'd333877839;
array[18380]=30'd557205073;
array[18381]=30'd406210138;
array[18382]=30'd406210138;
array[18383]=30'd417795660;
array[18384]=30'd641176139;
array[18385]=30'd883367490;
array[18386]=30'd959930934;
array[18387]=30'd959930934;
array[18388]=30'd959930934;
array[18389]=30'd641176139;
array[18390]=30'd597116464;
array[18391]=30'd548890196;
array[18392]=30'd548890196;
array[18393]=30'd548890196;
array[18394]=30'd571952708;
array[18395]=30'd548890196;
array[18396]=30'd548890196;
array[18397]=30'd548890196;
array[18398]=30'd707208791;
array[18399]=30'd883367490;
array[18400]=30'd959930934;
array[18401]=30'd959930934;
array[18402]=30'd959930934;
array[18403]=30'd959930934;
array[18404]=30'd883367490;
array[18405]=30'd624350812;
array[18406]=30'd362168943;
array[18407]=30'd637892242;
array[18408]=30'd452327079;
array[18409]=30'd601183923;
array[18410]=30'd548775573;
array[18411]=30'd373711515;
array[18412]=30'd463850128;
array[18413]=30'd637892242;
array[18414]=30'd556097214;
array[18415]=30'd779516542;
array[18416]=30'd879170165;
array[18417]=30'd857217603;
array[18418]=30'd820526616;
array[18419]=30'd809003452;
array[18420]=30'd965227994;
array[18421]=30'd983041534;
array[18422]=30'd894969309;
array[18423]=30'd785935846;
array[18424]=30'd767069629;
array[18425]=30'd767069629;
array[18426]=30'd767069629;
array[18427]=30'd792195525;
array[18428]=30'd871846383;
array[18429]=30'd883367490;
array[18430]=30'd879170165;
array[18431]=30'd879170165;
array[18432]=30'd900141674;
array[18433]=30'd900141674;
array[18434]=30'd900141674;
array[18435]=30'd900141674;
array[18436]=30'd900141674;
array[18437]=30'd900141674;
array[18438]=30'd900141674;
array[18439]=30'd900141674;
array[18440]=30'd879170165;
array[18441]=30'd879170165;
array[18442]=30'd900141674;
array[18443]=30'd900141674;
array[18444]=30'd900141674;
array[18445]=30'd900141674;
array[18446]=30'd900141674;
array[18447]=30'd900141674;
array[18448]=30'd804744750;
array[18449]=30'd409476630;
array[18450]=30'd492300766;
array[18451]=30'd475492838;
array[18452]=30'd804744750;
array[18453]=30'd900141674;
array[18454]=30'd900141674;
array[18455]=30'd900141674;
array[18456]=30'd900141674;
array[18457]=30'd900141674;
array[18458]=30'd900141674;
array[18459]=30'd900141674;
array[18460]=30'd900141674;
array[18461]=30'd824630873;
array[18462]=30'd468145703;
array[18463]=30'd492300766;
array[18464]=30'd490193319;
array[18465]=30'd490193319;
array[18466]=30'd448250284;
array[18467]=30'd414702010;
array[18468]=30'd414702010;
array[18469]=30'd448250284;
array[18470]=30'd461875644;
array[18471]=30'd461875644;
array[18472]=30'd394764738;
array[18473]=30'd359126474;
array[18474]=30'd422024669;
array[18475]=30'd422024669;
array[18476]=30'd422024669;
array[18477]=30'd371683842;
array[18478]=30'd300376570;
array[18479]=30'd333946399;
array[18480]=30'd333877839;
array[18481]=30'd449215039;
array[18482]=30'd679961142;
array[18483]=30'd916919852;
array[18484]=30'd959930934;
array[18485]=30'd859252262;
array[18486]=30'd804744750;
array[18487]=30'd941029952;
array[18488]=30'd883367490;
array[18489]=30'd859252262;
array[18490]=30'd859252262;
array[18491]=30'd842497613;
array[18492]=30'd916919852;
array[18493]=30'd959930934;
array[18494]=30'd959930934;
array[18495]=30'd959930934;
array[18496]=30'd959930934;
array[18497]=30'd959930934;
array[18498]=30'd916919852;
array[18499]=30'd751243845;
array[18500]=30'd449215039;
array[18501]=30'd406210138;
array[18502]=30'd446038641;
array[18503]=30'd583395966;
array[18504]=30'd518350503;
array[18505]=30'd601183923;
array[18506]=30'd427157133;
array[18507]=30'd322308749;
array[18508]=30'd463850128;
array[18509]=30'd637892242;
array[18510]=30'd548775573;
array[18511]=30'd855016073;
array[18512]=30'd879170165;
array[18513]=30'd900141674;
array[18514]=30'd857217603;
array[18515]=30'd785935846;
array[18516]=30'd832062938;
array[18517]=30'd965227994;
array[18518]=30'd983041534;
array[18519]=30'd916977147;
array[18520]=30'd872938009;
array[18521]=30'd855121400;
array[18522]=30'd855121400;
array[18523]=30'd893852174;
array[18524]=30'd916919852;
array[18525]=30'd883367490;
array[18526]=30'd879170165;
array[18527]=30'd879170165;
array[18528]=30'd900141674;
array[18529]=30'd900141674;
array[18530]=30'd900141674;
array[18531]=30'd900141674;
array[18532]=30'd900141674;
array[18533]=30'd900141674;
array[18534]=30'd900141674;
array[18535]=30'd900141674;
array[18536]=30'd900141674;
array[18537]=30'd900141674;
array[18538]=30'd900141674;
array[18539]=30'd900141674;
array[18540]=30'd900141674;
array[18541]=30'd900141674;
array[18542]=30'd900141674;
array[18543]=30'd900141674;
array[18544]=30'd842497613;
array[18545]=30'd517468675;
array[18546]=30'd777516526;
array[18547]=30'd839346691;
array[18548]=30'd792119862;
array[18549]=30'd900141674;
array[18550]=30'd900141674;
array[18551]=30'd900141674;
array[18552]=30'd900141674;
array[18553]=30'd900141674;
array[18554]=30'd900141674;
array[18555]=30'd900141674;
array[18556]=30'd883367490;
array[18557]=30'd571952708;
array[18558]=30'd492300766;
array[18559]=30'd479712691;
array[18560]=30'd490193319;
array[18561]=30'd490193319;
array[18562]=30'd490193319;
array[18563]=30'd490193319;
array[18564]=30'd479712691;
array[18565]=30'd479712691;
array[18566]=30'd479712691;
array[18567]=30'd479712691;
array[18568]=30'd461875644;
array[18569]=30'd372750770;
array[18570]=30'd479712691;
array[18571]=30'd479712691;
array[18572]=30'd461875644;
array[18573]=30'd461875644;
array[18574]=30'd394764738;
array[18575]=30'd422024669;
array[18576]=30'd316071465;
array[18577]=30'd449215039;
array[18578]=30'd406210138;
array[18579]=30'd417795660;
array[18580]=30'd571952708;
array[18581]=30'd722945572;
array[18582]=30'd665233987;
array[18583]=30'd941029952;
array[18584]=30'd959930934;
array[18585]=30'd959930934;
array[18586]=30'd959930934;
array[18587]=30'd979844654;
array[18588]=30'd959930934;
array[18589]=30'd979844654;
array[18590]=30'd959930934;
array[18591]=30'd941029952;
array[18592]=30'd883367490;
array[18593]=30'd792119862;
array[18594]=30'd510044739;
array[18595]=30'd449215039;
array[18596]=30'd446038641;
array[18597]=30'd406210138;
array[18598]=30'd503735925;
array[18599]=30'd463850128;
array[18600]=30'd611709603;
array[18601]=30'd497425057;
array[18602]=30'd322308749;
array[18603]=30'd289797789;
array[18604]=30'd503735925;
array[18605]=30'd637892242;
array[18606]=30'd559303301;
array[18607]=30'd879170165;
array[18608]=30'd879170165;
array[18609]=30'd879170165;
array[18610]=30'd898098744;
array[18611]=30'd857217603;
array[18612]=30'd785935846;
array[18613]=30'd832062938;
array[18614]=30'd965227994;
array[18615]=30'd983041534;
array[18616]=30'd936883742;
array[18617]=30'd936883742;
array[18618]=30'd936883742;
array[18619]=30'd959930934;
array[18620]=30'd941029952;
array[18621]=30'd879170165;
array[18622]=30'd879170165;
array[18623]=30'd900141674;
array[18624]=30'd900141674;
array[18625]=30'd900141674;
array[18626]=30'd900141674;
array[18627]=30'd900141674;
array[18628]=30'd900141674;
array[18629]=30'd900141674;
array[18630]=30'd900141674;
array[18631]=30'd900141674;
array[18632]=30'd900141674;
array[18633]=30'd900141674;
array[18634]=30'd900141674;
array[18635]=30'd900141674;
array[18636]=30'd900141674;
array[18637]=30'd900141674;
array[18638]=30'd900141674;
array[18639]=30'd900141674;
array[18640]=30'd857217603;
array[18641]=30'd737670674;
array[18642]=30'd1037554180;
array[18643]=30'd960978443;
array[18644]=30'd751243845;
array[18645]=30'd900141674;
array[18646]=30'd900141674;
array[18647]=30'd900141674;
array[18648]=30'd900141674;
array[18649]=30'd900141674;
array[18650]=30'd900141674;
array[18651]=30'd900141674;
array[18652]=30'd722945572;
array[18653]=30'd461903352;
array[18654]=30'd479712691;
array[18655]=30'd479712691;
array[18656]=30'd479712691;
array[18657]=30'd490193319;
array[18658]=30'd490193319;
array[18659]=30'd490193319;
array[18660]=30'd490193319;
array[18661]=30'd490193319;
array[18662]=30'd479712691;
array[18663]=30'd479712691;
array[18664]=30'd448250284;
array[18665]=30'd323471799;
array[18666]=30'd359126474;
array[18667]=30'd394764738;
array[18668]=30'd394764738;
array[18669]=30'd414702010;
array[18670]=30'd341278169;
array[18671]=30'd300376570;
array[18672]=30'd333877839;
array[18673]=30'd457612903;
array[18674]=30'd409377416;
array[18675]=30'd362168943;
array[18676]=30'd457612903;
array[18677]=30'd406210138;
array[18678]=30'd333877839;
array[18679]=30'd484882002;
array[18680]=30'd665233987;
array[18681]=30'd792119862;
array[18682]=30'd859252262;
array[18683]=30'd883367490;
array[18684]=30'd859252262;
array[18685]=30'd792119862;
array[18686]=30'd707208791;
array[18687]=30'd665233987;
array[18688]=30'd679961142;
array[18689]=30'd751243845;
array[18690]=30'd352806463;
array[18691]=30'd449215039;
array[18692]=30'd446038641;
array[18693]=30'd362168943;
array[18694]=30'd523632283;
array[18695]=30'd497425057;
array[18696]=30'd556097214;
array[18697]=30'd373711515;
array[18698]=30'd289797789;
array[18699]=30'd322308749;
array[18700]=30'd523632283;
array[18701]=30'd637892242;
array[18702]=30'd583395966;
array[18703]=30'd879170165;
array[18704]=30'd879170165;
array[18705]=30'd879170165;
array[18706]=30'd900141674;
array[18707]=30'd922198619;
array[18708]=30'd872938009;
array[18709]=30'd785935846;
array[18710]=30'd832062938;
array[18711]=30'd945318330;
array[18712]=30'd894969309;
array[18713]=30'd871910847;
array[18714]=30'd832062938;
array[18715]=30'd893852174;
array[18716]=30'd916919852;
array[18717]=30'd879170165;
array[18718]=30'd879170165;
array[18719]=30'd879170165;
array[18720]=30'd900141674;
array[18721]=30'd900141674;
array[18722]=30'd900141674;
array[18723]=30'd900141674;
array[18724]=30'd900141674;
array[18725]=30'd900141674;
array[18726]=30'd900141674;
array[18727]=30'd898098744;
array[18728]=30'd872938009;
array[18729]=30'd820526616;
array[18730]=30'd872938009;
array[18731]=30'd898098744;
array[18732]=30'd883367490;
array[18733]=30'd883367490;
array[18734]=30'd900141674;
array[18735]=30'd900141674;
array[18736]=30'd857217603;
array[18737]=30'd737670674;
array[18738]=30'd1037554180;
array[18739]=30'd996656669;
array[18740]=30'd751243845;
array[18741]=30'd900141674;
array[18742]=30'd900141674;
array[18743]=30'd900141674;
array[18744]=30'd900141674;
array[18745]=30'd900141674;
array[18746]=30'd900141674;
array[18747]=30'd842497613;
array[18748]=30'd461903352;
array[18749]=30'd492300766;
array[18750]=30'd479712691;
array[18751]=30'd479712691;
array[18752]=30'd414702010;
array[18753]=30'd448250284;
array[18754]=30'd448250284;
array[18755]=30'd461875644;
array[18756]=30'd479712691;
array[18757]=30'd490193319;
array[18758]=30'd479712691;
array[18759]=30'd490193319;
array[18760]=30'd479712691;
array[18761]=30'd461875644;
array[18762]=30'd359126474;
array[18763]=30'd414702010;
array[18764]=30'd394764738;
array[18765]=30'd300376570;
array[18766]=30'd378982955;
array[18767]=30'd248962651;
array[18768]=30'd406210138;
array[18769]=30'd433488509;
array[18770]=30'd409377416;
array[18771]=30'd362168943;
array[18772]=30'd446038641;
array[18773]=30'd433488509;
array[18774]=30'd409377416;
array[18775]=30'd337060463;
array[18776]=30'd406210138;
array[18777]=30'd484882002;
array[18778]=30'd792119862;
array[18779]=30'd792119862;
array[18780]=30'd792119862;
array[18781]=30'd792119862;
array[18782]=30'd794239590;
array[18783]=30'd824630873;
array[18784]=30'd824630873;
array[18785]=30'd751243845;
array[18786]=30'd237510232;
array[18787]=30'd314020436;
array[18788]=30'd406210138;
array[18789]=30'd433488509;
array[18790]=30'd463850128;
array[18791]=30'd611709603;
array[18792]=30'd444947126;
array[18793]=30'd337060463;
array[18794]=30'd373711515;
array[18795]=30'd362168943;
array[18796]=30'd523632283;
array[18797]=30'd601183923;
array[18798]=30'd651585154;
array[18799]=30'd879170165;
array[18800]=30'd900141674;
array[18801]=30'd879170165;
array[18802]=30'd879170165;
array[18803]=30'd900141674;
array[18804]=30'd898098744;
array[18805]=30'd872938009;
array[18806]=30'd785935846;
array[18807]=30'd753420739;
array[18808]=30'd767069629;
array[18809]=30'd792195525;
array[18810]=30'd815247846;
array[18811]=30'd893852174;
array[18812]=30'd883367490;
array[18813]=30'd900141674;
array[18814]=30'd879170165;
array[18815]=30'd879170165;
array[18816]=30'd900141674;
array[18817]=30'd900141674;
array[18818]=30'd900141674;
array[18819]=30'd900141674;
array[18820]=30'd900141674;
array[18821]=30'd900141674;
array[18822]=30'd898098744;
array[18823]=30'd820526616;
array[18824]=30'd832062938;
array[18825]=30'd832062938;
array[18826]=30'd809003452;
array[18827]=30'd785935846;
array[18828]=30'd815247846;
array[18829]=30'd872938009;
array[18830]=30'd883367490;
array[18831]=30'd900141674;
array[18832]=30'd898098744;
array[18833]=30'd650619404;
array[18834]=30'd1037554180;
array[18835]=30'd1037554180;
array[18836]=30'd722945572;
array[18837]=30'd900141674;
array[18838]=30'd900141674;
array[18839]=30'd900141674;
array[18840]=30'd900141674;
array[18841]=30'd900141674;
array[18842]=30'd900141674;
array[18843]=30'd679961142;
array[18844]=30'd517468675;
array[18845]=30'd492300766;
array[18846]=30'd479712691;
array[18847]=30'd589828536;
array[18848]=30'd753420739;
array[18849]=30'd809003452;
array[18850]=30'd753420739;
array[18851]=30'd619182551;
array[18852]=30'd525848010;
array[18853]=30'd479712691;
array[18854]=30'd414702010;
array[18855]=30'd414702010;
array[18856]=30'd414702010;
array[18857]=30'd394764738;
array[18858]=30'd341278169;
array[18859]=30'd341278169;
array[18860]=30'd396849695;
array[18861]=30'd449215039;
array[18862]=30'd449215039;
array[18863]=30'd298227292;
array[18864]=30'd406210138;
array[18865]=30'd446038641;
array[18866]=30'd406210138;
array[18867]=30'd265721461;
array[18868]=30'd446038641;
array[18869]=30'd446038641;
array[18870]=30'd427157133;
array[18871]=30'd362168943;
array[18872]=30'd298227292;
array[18873]=30'd352806463;
array[18874]=30'd824630873;
array[18875]=30'd824630873;
array[18876]=30'd824630873;
array[18877]=30'd824630873;
array[18878]=30'd824630873;
array[18879]=30'd794239590;
array[18880]=30'd679961142;
array[18881]=30'd417795660;
array[18882]=30'd268964427;
array[18883]=30'd268964427;
array[18884]=30'd248962651;
array[18885]=30'd446038641;
array[18886]=30'd523632283;
array[18887]=30'd548775573;
array[18888]=30'd373711515;
array[18889]=30'd337060463;
array[18890]=30'd406210138;
array[18891]=30'd362168943;
array[18892]=30'd523632283;
array[18893]=30'd611709603;
array[18894]=30'd681987696;
array[18895]=30'd879170165;
array[18896]=30'd879170165;
array[18897]=30'd879170165;
array[18898]=30'd900141674;
array[18899]=30'd879170165;
array[18900]=30'd900141674;
array[18901]=30'd900141674;
array[18902]=30'd857217603;
array[18903]=30'd872938009;
array[18904]=30'd872938009;
array[18905]=30'd893852174;
array[18906]=30'd916919852;
array[18907]=30'd883367490;
array[18908]=30'd900141674;
array[18909]=30'd900141674;
array[18910]=30'd879170165;
array[18911]=30'd879170165;
array[18912]=30'd900141674;
array[18913]=30'd900141674;
array[18914]=30'd900141674;
array[18915]=30'd900141674;
array[18916]=30'd900141674;
array[18917]=30'd922198619;
array[18918]=30'd820526616;
array[18919]=30'd855121400;
array[18920]=30'd983041534;
array[18921]=30'd1016593896;
array[18922]=30'd1016593896;
array[18923]=30'd948416998;
array[18924]=30'd832062938;
array[18925]=30'd792195525;
array[18926]=30'd871846383;
array[18927]=30'd916919852;
array[18928]=30'd936883742;
array[18929]=30'd737670674;
array[18930]=30'd983041534;
array[18931]=30'd1037554180;
array[18932]=30'd804744750;
array[18933]=30'd883367490;
array[18934]=30'd900141674;
array[18935]=30'd900141674;
array[18936]=30'd900141674;
array[18937]=30'd900141674;
array[18938]=30'd842497613;
array[18939]=30'd768057919;
array[18940]=30'd855121400;
array[18941]=30'd589828536;
array[18942]=30'd479712691;
array[18943]=30'd809003452;
array[18944]=30'd945318330;
array[18945]=30'd965227994;
array[18946]=30'd894969309;
array[18947]=30'd832062938;
array[18948]=30'd785935846;
array[18949]=30'd832062938;
array[18950]=30'd871910847;
array[18951]=30'd809003452;
array[18952]=30'd916977147;
array[18953]=30'd839346691;
array[18954]=30'd555187752;
array[18955]=30'd406210138;
array[18956]=30'd559303301;
array[18957]=30'd446038641;
array[18958]=30'd362168943;
array[18959]=30'd298227292;
array[18960]=30'd362168943;
array[18961]=30'd446038641;
array[18962]=30'd409377416;
array[18963]=30'd248962651;
array[18964]=30'd446038641;
array[18965]=30'd446038641;
array[18966]=30'd427157133;
array[18967]=30'd337060463;
array[18968]=30'd237510232;
array[18969]=30'd314020436;
array[18970]=30'd751243845;
array[18971]=30'd824630873;
array[18972]=30'd824630873;
array[18973]=30'd794239590;
array[18974]=30'd707208791;
array[18975]=30'd439898691;
array[18976]=30'd268964427;
array[18977]=30'd245976655;
array[18978]=30'd272186951;
array[18979]=30'd268964427;
array[18980]=30'd333877839;
array[18981]=30'd446038641;
array[18982]=30'd548775573;
array[18983]=30'd427157133;
array[18984]=30'd247877272;
array[18985]=30'd406210138;
array[18986]=30'd362168943;
array[18987]=30'd406210138;
array[18988]=30'd463850128;
array[18989]=30'd583395966;
array[18990]=30'd730239616;
array[18991]=30'd900141674;
array[18992]=30'd879170165;
array[18993]=30'd879170165;
array[18994]=30'd879170165;
array[18995]=30'd879170165;
array[18996]=30'd879170165;
array[18997]=30'd879170165;
array[18998]=30'd900141674;
array[18999]=30'd900141674;
array[19000]=30'd900141674;
array[19001]=30'd900141674;
array[19002]=30'd900141674;
array[19003]=30'd900141674;
array[19004]=30'd900141674;
array[19005]=30'd879170165;
array[19006]=30'd879170165;
array[19007]=30'd879170165;
array[19008]=30'd900141674;
array[19009]=30'd900141674;
array[19010]=30'd900141674;
array[19011]=30'd900141674;
array[19012]=30'd900141674;
array[19013]=30'd922198619;
array[19014]=30'd872938009;
array[19015]=30'd983041534;
array[19016]=30'd916977147;
array[19017]=30'd916977147;
array[19018]=30'd916977147;
array[19019]=30'd983041534;
array[19020]=30'd983041534;
array[19021]=30'd928507337;
array[19022]=30'd815247846;
array[19023]=30'd871846383;
array[19024]=30'd936883742;
array[19025]=30'd804744750;
array[19026]=30'd916977147;
array[19027]=30'd1037554180;
array[19028]=30'd872938009;
array[19029]=30'd804744750;
array[19030]=30'd900141674;
array[19031]=30'd900141674;
array[19032]=30'd900141674;
array[19033]=30'd900141674;
array[19034]=30'd725089870;
array[19035]=30'd996656669;
array[19036]=30'd1016593896;
array[19037]=30'd792195525;
array[19038]=30'd661135811;
array[19039]=30'd945318330;
array[19040]=30'd965227994;
array[19041]=30'd832062938;
array[19042]=30'd832062938;
array[19043]=30'd871910847;
array[19044]=30'd894969309;
array[19045]=30'd809003452;
array[19046]=30'd908629408;
array[19047]=30'd849905057;
array[19048]=30'd948416998;
array[19049]=30'd893852174;
array[19050]=30'd597116464;
array[19051]=30'd484882002;
array[19052]=30'd503735925;
array[19053]=30'd409377416;
array[19054]=30'd337060463;
array[19055]=30'd333877839;
array[19056]=30'd337060463;
array[19057]=30'd446038641;
array[19058]=30'd409377416;
array[19059]=30'd248962651;
array[19060]=30'd446038641;
array[19061]=30'd446038641;
array[19062]=30'd385301087;
array[19063]=30'd288874080;
array[19064]=30'd268964427;
array[19065]=30'd409476630;
array[19066]=30'd707208791;
array[19067]=30'd824630873;
array[19068]=30'd794239590;
array[19069]=30'd593953387;
array[19070]=30'd288874080;
array[19071]=30'd245976655;
array[19072]=30'd297344576;
array[19073]=30'd297344576;
array[19074]=30'd272186951;
array[19075]=30'd245976655;
array[19076]=30'd333877839;
array[19077]=30'd548775573;
array[19078]=30'd463850128;
array[19079]=30'd373711515;
array[19080]=30'd265721461;
array[19081]=30'd457612903;
array[19082]=30'd298227292;
array[19083]=30'd406210138;
array[19084]=30'd463850128;
array[19085]=30'd523632283;
array[19086]=30'd779516542;
array[19087]=30'd900141674;
array[19088]=30'd879170165;
array[19089]=30'd879170165;
array[19090]=30'd879170165;
array[19091]=30'd900141674;
array[19092]=30'd900141674;
array[19093]=30'd900141674;
array[19094]=30'd900141674;
array[19095]=30'd879170165;
array[19096]=30'd900141674;
array[19097]=30'd900141674;
array[19098]=30'd900141674;
array[19099]=30'd900141674;
array[19100]=30'd900141674;
array[19101]=30'd879170165;
array[19102]=30'd900141674;
array[19103]=30'd900141674;
array[19104]=30'd900141674;
array[19105]=30'd900141674;
array[19106]=30'd900141674;
array[19107]=30'd900141674;
array[19108]=30'd900141674;
array[19109]=30'd922198619;
array[19110]=30'd936883742;
array[19111]=30'd855121400;
array[19112]=30'd785935846;
array[19113]=30'd785935846;
array[19114]=30'd785935846;
array[19115]=30'd855121400;
array[19116]=30'd948416998;
array[19117]=30'd983041534;
array[19118]=30'd855121400;
array[19119]=30'd815247846;
array[19120]=30'd872938009;
array[19121]=30'd777516526;
array[19122]=30'd839346691;
array[19123]=30'd1037554180;
array[19124]=30'd960978443;
array[19125]=30'd722945572;
array[19126]=30'd900141674;
array[19127]=30'd900141674;
array[19128]=30'd900141674;
array[19129]=30'd900141674;
array[19130]=30'd842497613;
array[19131]=30'd996656669;
array[19132]=30'd983041534;
array[19133]=30'd709383649;
array[19134]=30'd832062938;
array[19135]=30'd965227994;
array[19136]=30'd894969309;
array[19137]=30'd785935846;
array[19138]=30'd945318330;
array[19139]=30'd894969309;
array[19140]=30'd945318330;
array[19141]=30'd809003452;
array[19142]=30'd893925805;
array[19143]=30'd849905057;
array[19144]=30'd948416998;
array[19145]=30'd893852174;
array[19146]=30'd583428668;
array[19147]=30'd614845038;
array[19148]=30'd373711515;
array[19149]=30'd373711515;
array[19150]=30'd333877839;
array[19151]=30'd362168943;
array[19152]=30'd337060463;
array[19153]=30'd446038641;
array[19154]=30'd457612903;
array[19155]=30'd333877839;
array[19156]=30'd337060463;
array[19157]=30'd314020436;
array[19158]=30'd268964427;
array[19159]=30'd288874080;
array[19160]=30'd230199867;
array[19161]=30'd395880013;
array[19162]=30'd804744750;
array[19163]=30'd768057919;
array[19164]=30'd503833159;
array[19165]=30'd268964427;
array[19166]=30'd272186951;
array[19167]=30'd297344576;
array[19168]=30'd297344576;
array[19169]=30'd272186951;
array[19170]=30'd297344576;
array[19171]=30'd268964427;
array[19172]=30'd457612903;
array[19173]=30'd548775573;
array[19174]=30'd427157133;
array[19175]=30'd265721461;
array[19176]=30'd385301087;
array[19177]=30'd457612903;
array[19178]=30'd298227292;
array[19179]=30'd406210138;
array[19180]=30'd463850128;
array[19181]=30'd523632283;
array[19182]=30'd779516542;
array[19183]=30'd900141674;
array[19184]=30'd879170165;
array[19185]=30'd879170165;
array[19186]=30'd900141674;
array[19187]=30'd900141674;
array[19188]=30'd900141674;
array[19189]=30'd900141674;
array[19190]=30'd900141674;
array[19191]=30'd900141674;
array[19192]=30'd879170165;
array[19193]=30'd900141674;
array[19194]=30'd900141674;
array[19195]=30'd900141674;
array[19196]=30'd900141674;
array[19197]=30'd879170165;
array[19198]=30'd900141674;
array[19199]=30'd900141674;
array[19200]=30'd900141674;
array[19201]=30'd900141674;
array[19202]=30'd900141674;
array[19203]=30'd900141674;
array[19204]=30'd900141674;
array[19205]=30'd922198619;
array[19206]=30'd898098744;
array[19207]=30'd785935846;
array[19208]=30'd832062938;
array[19209]=30'd894969309;
array[19210]=30'd871910847;
array[19211]=30'd767069629;
array[19212]=30'd894969309;
array[19213]=30'd948416998;
array[19214]=30'd916977147;
array[19215]=30'd785935846;
array[19216]=30'd894969309;
array[19217]=30'd916977147;
array[19218]=30'd737670674;
array[19219]=30'd1037554180;
array[19220]=30'd1037554180;
array[19221]=30'd722945572;
array[19222]=30'd916919852;
array[19223]=30'd900141674;
array[19224]=30'd900141674;
array[19225]=30'd900141674;
array[19226]=30'd922198619;
array[19227]=30'd959930934;
array[19228]=30'd820526616;
array[19229]=30'd777516526;
array[19230]=30'd832062938;
array[19231]=30'd965227994;
array[19232]=30'd855121400;
array[19233]=30'd832062938;
array[19234]=30'd945318330;
array[19235]=30'd767069629;
array[19236]=30'd792242589;
array[19237]=30'd829990281;
array[19238]=30'd849905057;
array[19239]=30'd871910847;
array[19240]=30'd948416998;
array[19241]=30'd916919852;
array[19242]=30'd557205073;
array[19243]=30'd637892242;
array[19244]=30'd373711515;
array[19245]=30'd362168943;
array[19246]=30'd298227292;
array[19247]=30'd406210138;
array[19248]=30'd337060463;
array[19249]=30'd337060463;
array[19250]=30'd352806463;
array[19251]=30'd268964427;
array[19252]=30'd237510232;
array[19253]=30'd230199867;
array[19254]=30'd241771065;
array[19255]=30'd272186951;
array[19256]=30'd241771065;
array[19257]=30'd268964427;
array[19258]=30'd725089870;
array[19259]=30'd439898691;
array[19260]=30'd241771065;
array[19261]=30'd272186951;
array[19262]=30'd272186951;
array[19263]=30'd272186951;
array[19264]=30'd272186951;
array[19265]=30'd272186951;
array[19266]=30'd241771065;
array[19267]=30'd298227292;
array[19268]=30'd559303301;
array[19269]=30'd463850128;
array[19270]=30'd362168943;
array[19271]=30'd223800938;
array[19272]=30'd298227292;
array[19273]=30'd337060463;
array[19274]=30'd298227292;
array[19275]=30'd362168943;
array[19276]=30'd463850128;
array[19277]=30'd523632283;
array[19278]=30'd824630873;
array[19279]=30'd900141674;
array[19280]=30'd879170165;
array[19281]=30'd879170165;
array[19282]=30'd900141674;
array[19283]=30'd900141674;
array[19284]=30'd900141674;
array[19285]=30'd900141674;
array[19286]=30'd900141674;
array[19287]=30'd900141674;
array[19288]=30'd879170165;
array[19289]=30'd900141674;
array[19290]=30'd900141674;
array[19291]=30'd900141674;
array[19292]=30'd900141674;
array[19293]=30'd900141674;
array[19294]=30'd900141674;
array[19295]=30'd900141674;
array[19296]=30'd900141674;
array[19297]=30'd900141674;
array[19298]=30'd900141674;
array[19299]=30'd900141674;
array[19300]=30'd900141674;
array[19301]=30'd900141674;
array[19302]=30'd898098744;
array[19303]=30'd820526616;
array[19304]=30'd965227994;
array[19305]=30'd945318330;
array[19306]=30'd945318330;
array[19307]=30'd871910847;
array[19308]=30'd809003452;
array[19309]=30'd894969309;
array[19310]=30'd916977147;
array[19311]=30'd785935846;
array[19312]=30'd894969309;
array[19313]=30'd983041534;
array[19314]=30'd709383649;
array[19315]=30'd1037554180;
array[19316]=30'd1037554180;
array[19317]=30'd804744750;
array[19318]=30'd883367490;
array[19319]=30'd900141674;
array[19320]=30'd900141674;
array[19321]=30'd900141674;
array[19322]=30'd900141674;
array[19323]=30'd883367490;
array[19324]=30'd725089870;
array[19325]=30'd898098744;
array[19326]=30'd820526616;
array[19327]=30'd916977147;
array[19328]=30'd894969309;
array[19329]=30'd832062938;
array[19330]=30'd945318330;
array[19331]=30'd849905057;
array[19332]=30'd908629408;
array[19333]=30'd849905057;
array[19334]=30'd871910847;
array[19335]=30'd948416998;
array[19336]=30'd916919852;
array[19337]=30'd883367490;
array[19338]=30'd557205073;
array[19339]=30'd637892242;
array[19340]=30'd427157133;
array[19341]=30'd265721461;
array[19342]=30'd298227292;
array[19343]=30'd352806463;
array[19344]=30'd395880013;
array[19345]=30'd453529185;
array[19346]=30'd439898691;
array[19347]=30'd346605135;
array[19348]=30'd272186951;
array[19349]=30'd241771065;
array[19350]=30'd297344576;
array[19351]=30'd297344576;
array[19352]=30'd272186951;
array[19353]=30'd206107200;
array[19354]=30'd327734842;
array[19355]=30'd268964427;
array[19356]=30'd272186951;
array[19357]=30'd297344576;
array[19358]=30'd272186951;
array[19359]=30'd272186951;
array[19360]=30'd272186951;
array[19361]=30'd272186951;
array[19362]=30'd268964427;
array[19363]=30'd484882002;
array[19364]=30'd503735925;
array[19365]=30'd427157133;
array[19366]=30'd337060463;
array[19367]=30'd248962651;
array[19368]=30'd268964427;
array[19369]=30'd268964427;
array[19370]=30'd218612285;
array[19371]=30'd333877839;
array[19372]=30'd446038641;
array[19373]=30'd497425057;
array[19374]=30'd794239590;
array[19375]=30'd900141674;
array[19376]=30'd879170165;
array[19377]=30'd879170165;
array[19378]=30'd900141674;
array[19379]=30'd900141674;
array[19380]=30'd900141674;
array[19381]=30'd900141674;
array[19382]=30'd900141674;
array[19383]=30'd900141674;
array[19384]=30'd900141674;
array[19385]=30'd900141674;
array[19386]=30'd900141674;
array[19387]=30'd900141674;
array[19388]=30'd900141674;
array[19389]=30'd900141674;
array[19390]=30'd879170165;
array[19391]=30'd900141674;
array[19392]=30'd900141674;
array[19393]=30'd900141674;
array[19394]=30'd900141674;
array[19395]=30'd900141674;
array[19396]=30'd900141674;
array[19397]=30'd900141674;
array[19398]=30'd898098744;
array[19399]=30'd820526616;
array[19400]=30'd871910847;
array[19401]=30'd792242589;
array[19402]=30'd871910847;
array[19403]=30'd945318330;
array[19404]=30'd809003452;
array[19405]=30'd809003452;
array[19406]=30'd965227994;
array[19407]=30'd785935846;
array[19408]=30'd832062938;
array[19409]=30'd855121400;
array[19410]=30'd666392059;
array[19411]=30'd948416998;
array[19412]=30'd1037554180;
array[19413]=30'd898098744;
array[19414]=30'd804744750;
array[19415]=30'd900141674;
array[19416]=30'd900141674;
array[19417]=30'd900141674;
array[19418]=30'd900141674;
array[19419]=30'd900141674;
array[19420]=30'd900141674;
array[19421]=30'd922198619;
array[19422]=30'd898098744;
array[19423]=30'd936883742;
array[19424]=30'd936883742;
array[19425]=30'd855121400;
array[19426]=30'd855121400;
array[19427]=30'd832062938;
array[19428]=30'd832062938;
array[19429]=30'd928507337;
array[19430]=30'd948416998;
array[19431]=30'd916919852;
array[19432]=30'd916919852;
array[19433]=30'd900141674;
array[19434]=30'd527849061;
array[19435]=30'd637892242;
array[19436]=30'd463850128;
array[19437]=30'd248962651;
array[19438]=30'd385301087;
array[19439]=30'd483946067;
array[19440]=30'd473528913;
array[19441]=30'd473528913;
array[19442]=30'd473528913;
array[19443]=30'd412708426;
array[19444]=30'd272186951;
array[19445]=30'd241771065;
array[19446]=30'd297344576;
array[19447]=30'd272186951;
array[19448]=30'd272186951;
array[19449]=30'd206107200;
array[19450]=30'd241771065;
array[19451]=30'd272186951;
array[19452]=30'd272186951;
array[19453]=30'd272186951;
array[19454]=30'd272186951;
array[19455]=30'd297344576;
array[19456]=30'd272186951;
array[19457]=30'd245976655;
array[19458]=30'd314020436;
array[19459]=30'd568787568;
array[19460]=30'd427157133;
array[19461]=30'd373711515;
array[19462]=30'd298227292;
array[19463]=30'd268964427;
array[19464]=30'd346605135;
array[19465]=30'd360280652;
array[19466]=30'd395880013;
array[19467]=30'd346605135;
array[19468]=30'd385301087;
array[19469]=30'd527849061;
array[19470]=30'd730239616;
array[19471]=30'd900141674;
array[19472]=30'd879170165;
array[19473]=30'd900141674;
array[19474]=30'd900141674;
array[19475]=30'd900141674;
array[19476]=30'd900141674;
array[19477]=30'd900141674;
array[19478]=30'd900141674;
array[19479]=30'd900141674;
array[19480]=30'd900141674;
array[19481]=30'd900141674;
array[19482]=30'd900141674;
array[19483]=30'd900141674;
array[19484]=30'd900141674;
array[19485]=30'd900141674;
array[19486]=30'd900141674;
array[19487]=30'd900141674;
array[19488]=30'd900141674;
array[19489]=30'd900141674;
array[19490]=30'd900141674;
array[19491]=30'd900141674;
array[19492]=30'd900141674;
array[19493]=30'd900141674;
array[19494]=30'd922198619;
array[19495]=30'd785935846;
array[19496]=30'd871910847;
array[19497]=30'd792242589;
array[19498]=30'd849905057;
array[19499]=30'd908629408;
array[19500]=30'd809003452;
array[19501]=30'd871910847;
array[19502]=30'd894969309;
array[19503]=30'd809003452;
array[19504]=30'd894969309;
array[19505]=30'd894969309;
array[19506]=30'd777516526;
array[19507]=30'd820526616;
array[19508]=30'd996656669;
array[19509]=30'd936883742;
array[19510]=30'd679961142;
array[19511]=30'd922198619;
array[19512]=30'd900141674;
array[19513]=30'd900141674;
array[19514]=30'd900141674;
array[19515]=30'd900141674;
array[19516]=30'd922198619;
array[19517]=30'd922198619;
array[19518]=30'd922198619;
array[19519]=30'd922198619;
array[19520]=30'd922198619;
array[19521]=30'd898098744;
array[19522]=30'd898098744;
array[19523]=30'd936883742;
array[19524]=30'd936883742;
array[19525]=30'd936883742;
array[19526]=30'd941029952;
array[19527]=30'd922198619;
array[19528]=30'd900141674;
array[19529]=30'd900141674;
array[19530]=30'd568787568;
array[19531]=30'd637892242;
array[19532]=30'd477520516;
array[19533]=30'd248962651;
array[19534]=30'd395880013;
array[19535]=30'd473528913;
array[19536]=30'd473528913;
array[19537]=30'd487155275;
array[19538]=30'd473528913;
array[19539]=30'd460936768;
array[19540]=30'd297344576;
array[19541]=30'd245976655;
array[19542]=30'd297344576;
array[19543]=30'd272186951;
array[19544]=30'd245976655;
array[19545]=30'd178845250;
array[19546]=30'd206107200;
array[19547]=30'd272186951;
array[19548]=30'd272186951;
array[19549]=30'd297344576;
array[19550]=30'd297344576;
array[19551]=30'd272186951;
array[19552]=30'd272186951;
array[19553]=30'd268964427;
array[19554]=30'd457612903;
array[19555]=30'd503735925;
array[19556]=30'd427157133;
array[19557]=30'd337060463;
array[19558]=30'd314020436;
array[19559]=30'd439898691;
array[19560]=30'd460936768;
array[19561]=30'd460936768;
array[19562]=30'd460936768;
array[19563]=30'd492371499;
array[19564]=30'd439898691;
array[19565]=30'd385301087;
array[19566]=30'd751243845;
array[19567]=30'd900141674;
array[19568]=30'd900141674;
array[19569]=30'd900141674;
array[19570]=30'd900141674;
array[19571]=30'd900141674;
array[19572]=30'd900141674;
array[19573]=30'd900141674;
array[19574]=30'd900141674;
array[19575]=30'd900141674;
array[19576]=30'd900141674;
array[19577]=30'd900141674;
array[19578]=30'd900141674;
array[19579]=30'd900141674;
array[19580]=30'd900141674;
array[19581]=30'd900141674;
array[19582]=30'd900141674;
array[19583]=30'd879170165;
array[19584]=30'd900141674;
array[19585]=30'd900141674;
array[19586]=30'd900141674;
array[19587]=30'd900141674;
array[19588]=30'd900141674;
array[19589]=30'd922198619;
array[19590]=30'd922198619;
array[19591]=30'd855121400;
array[19592]=30'd871910847;
array[19593]=30'd908629408;
array[19594]=30'd792242589;
array[19595]=30'd792242589;
array[19596]=30'd849905057;
array[19597]=30'd908629408;
array[19598]=30'd809003452;
array[19599]=30'd871910847;
array[19600]=30'd948416998;
array[19601]=30'd983041534;
array[19602]=30'd855121400;
array[19603]=30'd613923367;
array[19604]=30'd761730564;
array[19605]=30'd859252262;
array[19606]=30'd751243845;
array[19607]=30'd722945572;
array[19608]=30'd804744750;
array[19609]=30'd883367490;
array[19610]=30'd900141674;
array[19611]=30'd900141674;
array[19612]=30'd900141674;
array[19613]=30'd922198619;
array[19614]=30'd922198619;
array[19615]=30'd922198619;
array[19616]=30'd922198619;
array[19617]=30'd922198619;
array[19618]=30'd922198619;
array[19619]=30'd922198619;
array[19620]=30'd922198619;
array[19621]=30'd922198619;
array[19622]=30'd922198619;
array[19623]=30'd900141674;
array[19624]=30'd900141674;
array[19625]=30'd900141674;
array[19626]=30'd593953387;
array[19627]=30'd651585154;
array[19628]=30'd503735925;
array[19629]=30'd248962651;
array[19630]=30'd483946067;
array[19631]=30'd473528913;
array[19632]=30'd473528913;
array[19633]=30'd487155275;
array[19634]=30'd473528913;
array[19635]=30'd473528913;
array[19636]=30'd360280652;
array[19637]=30'd272186951;
array[19638]=30'd272186951;
array[19639]=30'd272186951;
array[19640]=30'd241771065;
array[19641]=30'd178845250;
array[19642]=30'd206107200;
array[19643]=30'd241771065;
array[19644]=30'd272186951;
array[19645]=30'd272186951;
array[19646]=30'd297344576;
array[19647]=30'd272186951;
array[19648]=30'd272186951;
array[19649]=30'd268964427;
array[19650]=30'd527849061;
array[19651]=30'd433488509;
array[19652]=30'd373711515;
array[19653]=30'd385301087;
array[19654]=30'd352806463;
array[19655]=30'd483946067;
array[19656]=30'd473528913;
array[19657]=30'd473528913;
array[19658]=30'd473528913;
array[19659]=30'd460936768;
array[19660]=30'd460936768;
array[19661]=30'd439898691;
array[19662]=30'd591943231;
array[19663]=30'd922198619;
array[19664]=30'd900141674;
array[19665]=30'd900141674;
array[19666]=30'd900141674;
array[19667]=30'd900141674;
array[19668]=30'd900141674;
array[19669]=30'd900141674;
array[19670]=30'd900141674;
array[19671]=30'd900141674;
array[19672]=30'd900141674;
array[19673]=30'd900141674;
array[19674]=30'd900141674;
array[19675]=30'd900141674;
array[19676]=30'd900141674;
array[19677]=30'd900141674;
array[19678]=30'd900141674;
array[19679]=30'd900141674;
array[19680]=30'd900141674;
array[19681]=30'd900141674;
array[19682]=30'd900141674;
array[19683]=30'd900141674;
array[19684]=30'd900141674;
array[19685]=30'd922198619;
array[19686]=30'd922198619;
array[19687]=30'd936883742;
array[19688]=30'd832062938;
array[19689]=30'd849905057;
array[19690]=30'd849905057;
array[19691]=30'd849905057;
array[19692]=30'd908629408;
array[19693]=30'd849905057;
array[19694]=30'd871910847;
array[19695]=30'd965227994;
array[19696]=30'd872938009;
array[19697]=30'd722945572;
array[19698]=30'd839346691;
array[19699]=30'd936883742;
array[19700]=30'd959930934;
array[19701]=30'd959930934;
array[19702]=30'd959930934;
array[19703]=30'd959930934;
array[19704]=30'd679961142;
array[19705]=30'd679961142;
array[19706]=30'd751243845;
array[19707]=30'd883367490;
array[19708]=30'd900141674;
array[19709]=30'd922198619;
array[19710]=30'd922198619;
array[19711]=30'd922198619;
array[19712]=30'd922198619;
array[19713]=30'd922198619;
array[19714]=30'd922198619;
array[19715]=30'd922198619;
array[19716]=30'd900141674;
array[19717]=30'd900141674;
array[19718]=30'd900141674;
array[19719]=30'd900141674;
array[19720]=30'd900141674;
array[19721]=30'd900141674;
array[19722]=30'd548890196;
array[19723]=30'd614845038;
array[19724]=30'd477520516;
array[19725]=30'd288874080;
array[19726]=30'd483946067;
array[19727]=30'd487155275;
array[19728]=30'd473528913;
array[19729]=30'd487155275;
array[19730]=30'd487155275;
array[19731]=30'd473528913;
array[19732]=30'd360280652;
array[19733]=30'd297344576;
array[19734]=30'd272186951;
array[19735]=30'd241771065;
array[19736]=30'd206107200;
array[19737]=30'd178845250;
array[19738]=30'd241771065;
array[19739]=30'd241771065;
array[19740]=30'd245976655;
array[19741]=30'd272186951;
array[19742]=30'd297344576;
array[19743]=30'd334045781;
array[19744]=30'd371776054;
array[19745]=30'd352806463;
array[19746]=30'd527849061;
array[19747]=30'd409377416;
array[19748]=30'd248962651;
array[19749]=30'd385301087;
array[19750]=30'd346605135;
array[19751]=30'd483946067;
array[19752]=30'd473528913;
array[19753]=30'd473528913;
array[19754]=30'd473528913;
array[19755]=30'd473528913;
array[19756]=30'd460936768;
array[19757]=30'd412708426;
array[19758]=30'd439898691;
array[19759]=30'd802671197;
array[19760]=30'd900141674;
array[19761]=30'd900141674;
array[19762]=30'd900141674;
array[19763]=30'd900141674;
array[19764]=30'd900141674;
array[19765]=30'd900141674;
array[19766]=30'd900141674;
array[19767]=30'd900141674;
array[19768]=30'd900141674;
array[19769]=30'd900141674;
array[19770]=30'd900141674;
array[19771]=30'd900141674;
array[19772]=30'd900141674;
array[19773]=30'd900141674;
array[19774]=30'd900141674;
array[19775]=30'd900141674;
array[19776]=30'd900141674;
array[19777]=30'd922198619;
array[19778]=30'd900141674;
array[19779]=30'd900141674;
array[19780]=30'd900141674;
array[19781]=30'd922198619;
array[19782]=30'd922198619;
array[19783]=30'd959930934;
array[19784]=30'd936883742;
array[19785]=30'd871910847;
array[19786]=30'd809003452;
array[19787]=30'd792242589;
array[19788]=30'd792242589;
array[19789]=30'd871910847;
array[19790]=30'd928507337;
array[19791]=30'd916977147;
array[19792]=30'd722945572;
array[19793]=30'd936883742;
array[19794]=30'd959930934;
array[19795]=30'd959930934;
array[19796]=30'd959930934;
array[19797]=30'd959930934;
array[19798]=30'd959930934;
array[19799]=30'd959930934;
array[19800]=30'd722945572;
array[19801]=30'd959930934;
array[19802]=30'd859252262;
array[19803]=30'd768057919;
array[19804]=30'd922198619;
array[19805]=30'd922198619;
array[19806]=30'd922198619;
array[19807]=30'd922198619;
array[19808]=30'd922198619;
array[19809]=30'd900141674;
array[19810]=30'd922198619;
array[19811]=30'd922198619;
array[19812]=30'd900141674;
array[19813]=30'd900141674;
array[19814]=30'd900141674;
array[19815]=30'd900141674;
array[19816]=30'd900141674;
array[19817]=30'd802671197;
array[19818]=30'd352806463;
array[19819]=30'd559303301;
array[19820]=30'd503735925;
array[19821]=30'd288874080;
array[19822]=30'd523825734;
array[19823]=30'd487155275;
array[19824]=30'd473528913;
array[19825]=30'd487155275;
array[19826]=30'd473528913;
array[19827]=30'd473528913;
array[19828]=30'd460936768;
array[19829]=30'd334045781;
array[19830]=30'd297344576;
array[19831]=30'd297344576;
array[19832]=30'd241771065;
array[19833]=30'd178845250;
array[19834]=30'd272186951;
array[19835]=30'd327734842;
array[19836]=30'd297344576;
array[19837]=30'd360280652;
array[19838]=30'd460936768;
array[19839]=30'd412708426;
array[19840]=30'd346605135;
array[19841]=30'd417795660;
array[19842]=30'd503735925;
array[19843]=30'd385301087;
array[19844]=30'd188150391;
array[19845]=30'd385301087;
array[19846]=30'd395880013;
array[19847]=30'd483946067;
array[19848]=30'd473528913;
array[19849]=30'd473528913;
array[19850]=30'd473528913;
array[19851]=30'd460936768;
array[19852]=30'd360280652;
array[19853]=30'd473528913;
array[19854]=30'd460936768;
array[19855]=30'd555256383;
array[19856]=30'd922198619;
array[19857]=30'd900141674;
array[19858]=30'd900141674;
array[19859]=30'd900141674;
array[19860]=30'd900141674;
array[19861]=30'd900141674;
array[19862]=30'd900141674;
array[19863]=30'd900141674;
array[19864]=30'd900141674;
array[19865]=30'd900141674;
array[19866]=30'd900141674;
array[19867]=30'd900141674;
array[19868]=30'd900141674;
array[19869]=30'd900141674;
array[19870]=30'd900141674;
array[19871]=30'd900141674;
array[19872]=30'd900141674;
array[19873]=30'd900141674;
array[19874]=30'd900141674;
array[19875]=30'd900141674;
array[19876]=30'd900141674;
array[19877]=30'd922198619;
array[19878]=30'd922198619;
array[19879]=30'd922198619;
array[19880]=30'd959930934;
array[19881]=30'd936883742;
array[19882]=30'd983041534;
array[19883]=30'd894969309;
array[19884]=30'd928507337;
array[19885]=30'd948416998;
array[19886]=30'd936883742;
array[19887]=30'd916919852;
array[19888]=30'd768057919;
array[19889]=30'd979844654;
array[19890]=30'd959930934;
array[19891]=30'd959930934;
array[19892]=30'd959930934;
array[19893]=30'd959930934;
array[19894]=30'd959930934;
array[19895]=30'd941029952;
array[19896]=30'd751243845;
array[19897]=30'd959930934;
array[19898]=30'd916919852;
array[19899]=30'd751243845;
array[19900]=30'd922198619;
array[19901]=30'd922198619;
array[19902]=30'd922198619;
array[19903]=30'd922198619;
array[19904]=30'd922198619;
array[19905]=30'd922198619;
array[19906]=30'd922198619;
array[19907]=30'd922198619;
array[19908]=30'd922198619;
array[19909]=30'd922198619;
array[19910]=30'd900141674;
array[19911]=30'd900141674;
array[19912]=30'd900141674;
array[19913]=30'd575153766;
array[19914]=30'd453529185;
array[19915]=30'd484882002;
array[19916]=30'd503735925;
array[19917]=30'd268964427;
array[19918]=30'd483946067;
array[19919]=30'd473528913;
array[19920]=30'd487155275;
array[19921]=30'd487155275;
array[19922]=30'd487155275;
array[19923]=30'd487155275;
array[19924]=30'd473528913;
array[19925]=30'd473528913;
array[19926]=30'd473528913;
array[19927]=30'd460936768;
array[19928]=30'd360280652;
array[19929]=30'd245976655;
array[19930]=30'd412708426;
array[19931]=30'd460936768;
array[19932]=30'd460936768;
array[19933]=30'd412708426;
array[19934]=30'd360280652;
array[19935]=30'd360280652;
array[19936]=30'd439898691;
array[19937]=30'd484882002;
array[19938]=30'd457612903;
array[19939]=30'd288874080;
array[19940]=30'd237510232;
array[19941]=30'd385301087;
array[19942]=30'd439898691;
array[19943]=30'd460936768;
array[19944]=30'd473528913;
array[19945]=30'd473528913;
array[19946]=30'd460936768;
array[19947]=30'd412708426;
array[19948]=30'd460936768;
array[19949]=30'd473528913;
array[19950]=30'd473528913;
array[19951]=30'd412708426;
array[19952]=30'd842497613;
array[19953]=30'd922198619;
array[19954]=30'd900141674;
array[19955]=30'd900141674;
array[19956]=30'd900141674;
array[19957]=30'd900141674;
array[19958]=30'd900141674;
array[19959]=30'd900141674;
array[19960]=30'd900141674;
array[19961]=30'd922198619;
array[19962]=30'd922198619;
array[19963]=30'd922198619;
array[19964]=30'd922198619;
array[19965]=30'd900141674;
array[19966]=30'd922198619;
array[19967]=30'd900141674;
array[19968]=30'd900141674;
array[19969]=30'd900141674;
array[19970]=30'd900141674;
array[19971]=30'd900141674;
array[19972]=30'd922198619;
array[19973]=30'd922198619;
array[19974]=30'd922198619;
array[19975]=30'd922198619;
array[19976]=30'd922198619;
array[19977]=30'd922198619;
array[19978]=30'd959930934;
array[19979]=30'd959930934;
array[19980]=30'd959930934;
array[19981]=30'd959930934;
array[19982]=30'd922198619;
array[19983]=30'd922198619;
array[19984]=30'd804744750;
array[19985]=30'd959930934;
array[19986]=30'd959930934;
array[19987]=30'd959930934;
array[19988]=30'd959930934;
array[19989]=30'd959930934;
array[19990]=30'd959930934;
array[19991]=30'd959930934;
array[19992]=30'd751243845;
array[19993]=30'd959930934;
array[19994]=30'd859252262;
array[19995]=30'd804744750;
array[19996]=30'd922198619;
array[19997]=30'd922198619;
array[19998]=30'd922198619;
array[19999]=30'd922198619;
array[20000]=30'd922198619;
array[20001]=30'd922198619;
array[20002]=30'd922198619;
array[20003]=30'd922198619;
array[20004]=30'd922198619;
array[20005]=30'd922198619;
array[20006]=30'd922198619;
array[20007]=30'd922198619;
array[20008]=30'd802671197;
array[20009]=30'd439898691;
array[20010]=30'd483946067;
array[20011]=30'd395880013;
array[20012]=30'd453529185;
array[20013]=30'd268964427;
array[20014]=30'd483946067;
array[20015]=30'd473528913;
array[20016]=30'd487155275;
array[20017]=30'd487155275;
array[20018]=30'd487155275;
array[20019]=30'd487155275;
array[20020]=30'd473528913;
array[20021]=30'd473528913;
array[20022]=30'd473528913;
array[20023]=30'd473528913;
array[20024]=30'd460936768;
array[20025]=30'd297344576;
array[20026]=30'd460936768;
array[20027]=30'd473528913;
array[20028]=30'd473528913;
array[20029]=30'd473528913;
array[20030]=30'd460936768;
array[20031]=30'd460936768;
array[20032]=30'd460936768;
array[20033]=30'd439898691;
array[20034]=30'd457612903;
array[20035]=30'd288874080;
array[20036]=30'd395880013;
array[20037]=30'd288874080;
array[20038]=30'd439898691;
array[20039]=30'd473528913;
array[20040]=30'd473528913;
array[20041]=30'd473528913;
array[20042]=30'd412708426;
array[20043]=30'd460936768;
array[20044]=30'd473528913;
array[20045]=30'd473528913;
array[20046]=30'd473528913;
array[20047]=30'd460936768;
array[20048]=30'd697839152;
array[20049]=30'd922198619;
array[20050]=30'd900141674;
array[20051]=30'd900141674;
array[20052]=30'd900141674;
array[20053]=30'd922198619;
array[20054]=30'd900141674;
array[20055]=30'd922198619;
array[20056]=30'd922198619;
array[20057]=30'd922198619;
array[20058]=30'd959930934;
array[20059]=30'd936883742;
array[20060]=30'd872938009;
array[20061]=30'd872938009;
array[20062]=30'd872938009;
array[20063]=30'd898098744;
array[20064]=30'd922198619;
array[20065]=30'd900141674;
array[20066]=30'd922198619;
array[20067]=30'd922198619;
array[20068]=30'd922198619;
array[20069]=30'd922198619;
array[20070]=30'd922198619;
array[20071]=30'd922198619;
array[20072]=30'd922198619;
array[20073]=30'd922198619;
array[20074]=30'd922198619;
array[20075]=30'd922198619;
array[20076]=30'd922198619;
array[20077]=30'd922198619;
array[20078]=30'd922198619;
array[20079]=30'd900141674;
array[20080]=30'd768057919;
array[20081]=30'd959930934;
array[20082]=30'd959930934;
array[20083]=30'd979844654;
array[20084]=30'd959930934;
array[20085]=30'd959930934;
array[20086]=30'd959930934;
array[20087]=30'd959930934;
array[20088]=30'd768057919;
array[20089]=30'd804744750;
array[20090]=30'd641176139;
array[20091]=30'd883367490;
array[20092]=30'd922198619;
array[20093]=30'd922198619;
array[20094]=30'd922198619;
array[20095]=30'd922198619;
array[20096]=30'd922198619;
array[20097]=30'd922198619;
array[20098]=30'd922198619;
array[20099]=30'd922198619;
array[20100]=30'd922198619;
array[20101]=30'd922198619;
array[20102]=30'd922198619;
array[20103]=30'd883367490;
array[20104]=30'd521646692;
array[20105]=30'd460936768;
array[20106]=30'd473528913;
array[20107]=30'd483946067;
array[20108]=30'd346605135;
array[20109]=30'd268964427;
array[20110]=30'd395880013;
array[20111]=30'd473528913;
array[20112]=30'd487155275;
array[20113]=30'd487155275;
array[20114]=30'd487155275;
array[20115]=30'd487155275;
array[20116]=30'd487155275;
array[20117]=30'd473528913;
array[20118]=30'd473528913;
array[20119]=30'd473528913;
array[20120]=30'd360280652;
array[20121]=30'd334045781;
array[20122]=30'd473528913;
array[20123]=30'd473528913;
array[20124]=30'd473528913;
array[20125]=30'd473528913;
array[20126]=30'd473528913;
array[20127]=30'd473528913;
array[20128]=30'd460936768;
array[20129]=30'd346605135;
array[20130]=30'd352806463;
array[20131]=30'd395880013;
array[20132]=30'd483946067;
array[20133]=30'd346605135;
array[20134]=30'd395880013;
array[20135]=30'd473528913;
array[20136]=30'd473528913;
array[20137]=30'd460936768;
array[20138]=30'd412708426;
array[20139]=30'd473528913;
array[20140]=30'd473528913;
array[20141]=30'd473528913;
array[20142]=30'd473528913;
array[20143]=30'd460936768;
array[20144]=30'd591943231;
array[20145]=30'd922198619;
array[20146]=30'd900141674;
array[20147]=30'd900141674;
array[20148]=30'd900141674;
array[20149]=30'd922198619;
array[20150]=30'd922198619;
array[20151]=30'd922198619;
array[20152]=30'd979844654;
array[20153]=30'd936883742;
array[20154]=30'd809003452;
array[20155]=30'd767069629;
array[20156]=30'd778590630;
array[20157]=30'd778590630;
array[20158]=30'd767069629;
array[20159]=30'd767069629;
array[20160]=30'd941029952;
array[20161]=30'd922198619;
array[20162]=30'd922198619;
array[20163]=30'd922198619;
array[20164]=30'd922198619;
array[20165]=30'd922198619;
array[20166]=30'd922198619;
array[20167]=30'd922198619;
array[20168]=30'd922198619;
array[20169]=30'd922198619;
array[20170]=30'd922198619;
array[20171]=30'd922198619;
array[20172]=30'd900141674;
array[20173]=30'd922198619;
array[20174]=30'd922198619;
array[20175]=30'd922198619;
array[20176]=30'd707208791;
array[20177]=30'd959930934;
array[20178]=30'd959930934;
array[20179]=30'd979844654;
array[20180]=30'd979844654;
array[20181]=30'd959930934;
array[20182]=30'd959930934;
array[20183]=30'd959930934;
array[20184]=30'd959930934;
array[20185]=30'd842497613;
array[20186]=30'd883367490;
array[20187]=30'd922198619;
array[20188]=30'd922198619;
array[20189]=30'd922198619;
array[20190]=30'd922198619;
array[20191]=30'd922198619;
array[20192]=30'd922198619;
array[20193]=30'd922198619;
array[20194]=30'd922198619;
array[20195]=30'd922198619;
array[20196]=30'd922198619;
array[20197]=30'd922198619;
array[20198]=30'd898098744;
array[20199]=30'd503833159;
array[20200]=30'd483946067;
array[20201]=30'd473528913;
array[20202]=30'd487155275;
array[20203]=30'd487155275;
array[20204]=30'd395880013;
array[20205]=30'd268964427;
array[20206]=30'd439898691;
array[20207]=30'd473528913;
array[20208]=30'd487155275;
array[20209]=30'd487155275;
array[20210]=30'd487155275;
array[20211]=30'd487155275;
array[20212]=30'd473528913;
array[20213]=30'd473528913;
array[20214]=30'd473528913;
array[20215]=30'd460936768;
array[20216]=30'd360280652;
array[20217]=30'd360280652;
array[20218]=30'd473528913;
array[20219]=30'd473528913;
array[20220]=30'd473528913;
array[20221]=30'd473528913;
array[20222]=30'd487155275;
array[20223]=30'd473528913;
array[20224]=30'd473528913;
array[20225]=30'd371776054;
array[20226]=30'd288874080;
array[20227]=30'd483946067;
array[20228]=30'd460936768;
array[20229]=30'd460936768;
array[20230]=30'd334045781;
array[20231]=30'd460936768;
array[20232]=30'd473528913;
array[20233]=30'd360280652;
array[20234]=30'd473528913;
array[20235]=30'd473528913;
array[20236]=30'd473528913;
array[20237]=30'd473528913;
array[20238]=30'd473528913;
array[20239]=30'd473528913;
array[20240]=30'd483946067;
array[20241]=30'd898098744;
array[20242]=30'd922198619;
array[20243]=30'd922198619;
array[20244]=30'd922198619;
array[20245]=30'd922198619;
array[20246]=30'd922198619;
array[20247]=30'd979844654;
array[20248]=30'd936883742;
array[20249]=30'd809003452;
array[20250]=30'd792242589;
array[20251]=30'd829990281;
array[20252]=30'd849905057;
array[20253]=30'd849905057;
array[20254]=30'd908629408;
array[20255]=30'd849905057;
array[20256]=30'd916977147;
array[20257]=30'd936883742;
array[20258]=30'd922198619;
array[20259]=30'd922198619;
array[20260]=30'd922198619;
array[20261]=30'd922198619;
array[20262]=30'd922198619;
array[20263]=30'd922198619;
array[20264]=30'd922198619;
array[20265]=30'd922198619;
array[20266]=30'd922198619;
array[20267]=30'd922198619;
array[20268]=30'd922198619;
array[20269]=30'd922198619;
array[20270]=30'd922198619;
array[20271]=30'd922198619;
array[20272]=30'd725089870;
array[20273]=30'd959930934;
array[20274]=30'd979844654;
array[20275]=30'd979844654;
array[20276]=30'd979844654;
array[20277]=30'd959930934;
array[20278]=30'd959930934;
array[20279]=30'd959930934;
array[20280]=30'd959930934;
array[20281]=30'd804744750;
array[20282]=30'd883367490;
array[20283]=30'd922198619;
array[20284]=30'd922198619;
array[20285]=30'd922198619;
array[20286]=30'd922198619;
array[20287]=30'd922198619;
array[20288]=30'd922198619;
array[20289]=30'd922198619;
array[20290]=30'd922198619;
array[20291]=30'd922198619;
array[20292]=30'd922198619;
array[20293]=30'd922198619;
array[20294]=30'd591943231;
array[20295]=30'd460936768;
array[20296]=30'd487155275;
array[20297]=30'd487155275;
array[20298]=30'd487155275;
array[20299]=30'd487155275;
array[20300]=30'd412708426;
array[20301]=30'd327734842;
array[20302]=30'd395880013;
array[20303]=30'd473528913;
array[20304]=30'd487155275;
array[20305]=30'd487155275;
array[20306]=30'd487155275;
array[20307]=30'd487155275;
array[20308]=30'd487155275;
array[20309]=30'd473528913;
array[20310]=30'd473528913;
array[20311]=30'd360280652;
array[20312]=30'd412708426;
array[20313]=30'd360280652;
array[20314]=30'd473528913;
array[20315]=30'd473528913;
array[20316]=30'd473528913;
array[20317]=30'd473528913;
array[20318]=30'd487155275;
array[20319]=30'd487155275;
array[20320]=30'd473528913;
array[20321]=30'd412708426;
array[20322]=30'd241771065;
array[20323]=30'd460936768;
array[20324]=30'd473528913;
array[20325]=30'd473528913;
array[20326]=30'd460936768;
array[20327]=30'd460936768;
array[20328]=30'd412708426;
array[20329]=30'd412708426;
array[20330]=30'd473528913;
array[20331]=30'd473528913;
array[20332]=30'd473528913;
array[20333]=30'd473528913;
array[20334]=30'd473528913;
array[20335]=30'd473528913;
array[20336]=30'd412708426;
array[20337]=30'd842497613;
array[20338]=30'd922198619;
array[20339]=30'd922198619;
array[20340]=30'd922198619;
array[20341]=30'd922198619;
array[20342]=30'd959930934;
array[20343]=30'd983041534;
array[20344]=30'd832062938;
array[20345]=30'd792242589;
array[20346]=30'd908629408;
array[20347]=30'd908629408;
array[20348]=30'd792242589;
array[20349]=30'd792242589;
array[20350]=30'd945318330;
array[20351]=30'd945318330;
array[20352]=30'd871910847;
array[20353]=30'd916977147;
array[20354]=30'd941029952;
array[20355]=30'd922198619;
array[20356]=30'd922198619;
array[20357]=30'd922198619;
array[20358]=30'd922198619;
array[20359]=30'd922198619;
array[20360]=30'd922198619;
array[20361]=30'd922198619;
array[20362]=30'd922198619;
array[20363]=30'd922198619;
array[20364]=30'd922198619;
array[20365]=30'd922198619;
array[20366]=30'd922198619;
array[20367]=30'd922198619;
array[20368]=30'd768057919;
array[20369]=30'd898098744;
array[20370]=30'd959930934;
array[20371]=30'd959930934;
array[20372]=30'd979844654;
array[20373]=30'd959930934;
array[20374]=30'd959930934;
array[20375]=30'd979844654;
array[20376]=30'd959930934;
array[20377]=30'd722945572;
array[20378]=30'd722945572;
array[20379]=30'd941029952;
array[20380]=30'd922198619;
array[20381]=30'd922198619;
array[20382]=30'd922198619;
array[20383]=30'd922198619;
array[20384]=30'd922198619;
array[20385]=30'd922198619;
array[20386]=30'd922198619;
array[20387]=30'd922198619;
array[20388]=30'd922198619;
array[20389]=30'd609756759;
array[20390]=30'd460936768;
array[20391]=30'd487155275;
array[20392]=30'd487155275;
array[20393]=30'd487155275;
array[20394]=30'd473528913;
array[20395]=30'd460936768;
array[20396]=30'd412708426;
array[20397]=30'd460936768;
array[20398]=30'd360280652;
array[20399]=30'd460936768;
array[20400]=30'd473528913;
array[20401]=30'd487155275;
array[20402]=30'd487155275;
array[20403]=30'd487155275;
array[20404]=30'd473528913;
array[20405]=30'd473528913;
array[20406]=30'd460936768;
array[20407]=30'd360280652;
array[20408]=30'd460936768;
array[20409]=30'd412708426;
array[20410]=30'd473528913;
array[20411]=30'd473528913;
array[20412]=30'd473528913;
array[20413]=30'd473528913;
array[20414]=30'd487155275;
array[20415]=30'd473528913;
array[20416]=30'd460936768;
array[20417]=30'd483946067;
array[20418]=30'd327734842;
array[20419]=30'd483946067;
array[20420]=30'd487155275;
array[20421]=30'd473528913;
array[20422]=30'd473528913;
array[20423]=30'd460936768;
array[20424]=30'd360280652;
array[20425]=30'd460936768;
array[20426]=30'd473528913;
array[20427]=30'd473528913;
array[20428]=30'd473528913;
array[20429]=30'd473528913;
array[20430]=30'd473528913;
array[20431]=30'd473528913;
array[20432]=30'd412708426;
array[20433]=30'd725089870;
array[20434]=30'd922198619;
array[20435]=30'd922198619;
array[20436]=30'd922198619;
array[20437]=30'd959930934;
array[20438]=30'd996656669;
array[20439]=30'd832062938;
array[20440]=30'd792242589;
array[20441]=30'd876132737;
array[20442]=30'd829990281;
array[20443]=30'd766030218;
array[20444]=30'd766030218;
array[20445]=30'd766030218;
array[20446]=30'd871910847;
array[20447]=30'd997736898;
array[20448]=30'd809003452;
array[20449]=30'd832062938;
array[20450]=30'd936883742;
array[20451]=30'd941029952;
array[20452]=30'd922198619;
array[20453]=30'd922198619;
array[20454]=30'd922198619;
array[20455]=30'd922198619;
array[20456]=30'd922198619;
array[20457]=30'd922198619;
array[20458]=30'd922198619;
array[20459]=30'd922198619;
array[20460]=30'd922198619;
array[20461]=30'd922198619;
array[20462]=30'd922198619;
array[20463]=30'd922198619;
array[20464]=30'd857217603;
array[20465]=30'd804744750;
array[20466]=30'd959930934;
array[20467]=30'd959930934;
array[20468]=30'd959930934;
array[20469]=30'd959930934;
array[20470]=30'd959930934;
array[20471]=30'd959930934;
array[20472]=30'd959930934;
array[20473]=30'd679961142;
array[20474]=30'd768057919;
array[20475]=30'd859252262;
array[20476]=30'd922198619;
array[20477]=30'd922198619;
array[20478]=30'd922198619;
array[20479]=30'd922198619;
array[20480]=30'd922198619;
array[20481]=30'd922198619;
array[20482]=30'd922198619;
array[20483]=30'd922198619;
array[20484]=30'd609756759;
array[20485]=30'd483946067;
array[20486]=30'd487155275;
array[20487]=30'd487155275;
array[20488]=30'd473528913;
array[20489]=30'd473528913;
array[20490]=30'd460936768;
array[20491]=30'd412708426;
array[20492]=30'd473528913;
array[20493]=30'd473528913;
array[20494]=30'd473528913;
array[20495]=30'd460936768;
array[20496]=30'd473528913;
array[20497]=30'd487155275;
array[20498]=30'd487155275;
array[20499]=30'd487155275;
array[20500]=30'd473528913;
array[20501]=30'd473528913;
array[20502]=30'd360280652;
array[20503]=30'd460936768;
array[20504]=30'd412708426;
array[20505]=30'd412708426;
array[20506]=30'd473528913;
array[20507]=30'd473528913;
array[20508]=30'd473528913;
array[20509]=30'd473528913;
array[20510]=30'd487155275;
array[20511]=30'd473528913;
array[20512]=30'd555256383;
array[20513]=30'd842497613;
array[20514]=30'd641176139;
array[20515]=30'd656960070;
array[20516]=30'd483946067;
array[20517]=30'd460936768;
array[20518]=30'd473528913;
array[20519]=30'd460936768;
array[20520]=30'd334045781;
array[20521]=30'd460936768;
array[20522]=30'd412708426;
array[20523]=30'd460936768;
array[20524]=30'd473528913;
array[20525]=30'd473528913;
array[20526]=30'd473528913;
array[20527]=30'd487155275;
array[20528]=30'd473528913;
array[20529]=30'd483946067;
array[20530]=30'd898098744;
array[20531]=30'd922198619;
array[20532]=30'd922198619;
array[20533]=30'd979844654;
array[20534]=30'd916977147;
array[20535]=30'd767069629;
array[20536]=30'd829990281;
array[20537]=30'd829990281;
array[20538]=30'd766030218;
array[20539]=30'd829990281;
array[20540]=30'd908629408;
array[20541]=30'd849905057;
array[20542]=30'd893925805;
array[20543]=30'd977825191;
array[20544]=30'd945318330;
array[20545]=30'd809003452;
array[20546]=30'd894969309;
array[20547]=30'd936883742;
array[20548]=30'd941029952;
array[20549]=30'd922198619;
array[20550]=30'd922198619;
array[20551]=30'd922198619;
array[20552]=30'd922198619;
array[20553]=30'd922198619;
array[20554]=30'd922198619;
array[20555]=30'd922198619;
array[20556]=30'd922198619;
array[20557]=30'd922198619;
array[20558]=30'd922198619;
array[20559]=30'd922198619;
array[20560]=30'd922198619;
array[20561]=30'd768057919;
array[20562]=30'd898098744;
array[20563]=30'd959930934;
array[20564]=30'd959930934;
array[20565]=30'd959930934;
array[20566]=30'd959930934;
array[20567]=30'd959930934;
array[20568]=30'd859252262;
array[20569]=30'd804744750;
array[20570]=30'd959930934;
array[20571]=30'd768057919;
array[20572]=30'd883367490;
array[20573]=30'd922198619;
array[20574]=30'd922198619;
array[20575]=30'd922198619;
array[20576]=30'd922198619;
array[20577]=30'd922198619;
array[20578]=30'd922198619;
array[20579]=30'd725089870;
array[20580]=30'd439898691;
array[20581]=30'd492371499;
array[20582]=30'd487155275;
array[20583]=30'd487155275;
array[20584]=30'd487155275;
array[20585]=30'd460936768;
array[20586]=30'd412708426;
array[20587]=30'd473528913;
array[20588]=30'd473528913;
array[20589]=30'd487155275;
array[20590]=30'd487155275;
array[20591]=30'd487155275;
array[20592]=30'd473528913;
array[20593]=30'd487155275;
array[20594]=30'd487155275;
array[20595]=30'd473528913;
array[20596]=30'd360280652;
array[20597]=30'd412708426;
array[20598]=30'd360280652;
array[20599]=30'd473528913;
array[20600]=30'd412708426;
array[20601]=30'd460936768;
array[20602]=30'd473528913;
array[20603]=30'd473528913;
array[20604]=30'd473528913;
array[20605]=30'd487155275;
array[20606]=30'd473528913;
array[20607]=30'd523825734;
array[20608]=30'd842497613;
array[20609]=30'd597116464;
array[20610]=30'd679961142;
array[20611]=30'd641176139;
array[20612]=30'd483946067;
array[20613]=30'd460936768;
array[20614]=30'd460936768;
array[20615]=30'd422122009;
array[20616]=30'd820526616;
array[20617]=30'd936883742;
array[20618]=30'd898098744;
array[20619]=30'd555256383;
array[20620]=30'd460936768;
array[20621]=30'd473528913;
array[20622]=30'd487155275;
array[20623]=30'd473528913;
array[20624]=30'd473528913;
array[20625]=30'd460936768;
array[20626]=30'd725089870;
array[20627]=30'd936883742;
array[20628]=30'd959930934;
array[20629]=30'd979844654;
array[20630]=30'd916977147;
array[20631]=30'd767069629;
array[20632]=30'd876132737;
array[20633]=30'd792242589;
array[20634]=30'd766030218;
array[20635]=30'd908629408;
array[20636]=30'd977825191;
array[20637]=30'd997736898;
array[20638]=30'd908629408;
array[20639]=30'd809003452;
array[20640]=30'd945318330;
array[20641]=30'd792195525;
array[20642]=30'd894969309;
array[20643]=30'd983041534;
array[20644]=30'd872938009;
array[20645]=30'd941029952;
array[20646]=30'd922198619;
array[20647]=30'd922198619;
array[20648]=30'd922198619;
array[20649]=30'd922198619;
array[20650]=30'd922198619;
array[20651]=30'd922198619;
array[20652]=30'd922198619;
array[20653]=30'd922198619;
array[20654]=30'd922198619;
array[20655]=30'd922198619;
array[20656]=30'd922198619;
array[20657]=30'd900141674;
array[20658]=30'd768057919;
array[20659]=30'd916919852;
array[20660]=30'd959930934;
array[20661]=30'd959930934;
array[20662]=30'd936883742;
array[20663]=30'd804744750;
array[20664]=30'd722945572;
array[20665]=30'd959930934;
array[20666]=30'd959930934;
array[20667]=30'd959930934;
array[20668]=30'd768057919;
array[20669]=30'd922198619;
array[20670]=30'd922198619;
array[20671]=30'd922198619;
array[20672]=30'd922198619;
array[20673]=30'd922198619;
array[20674]=30'd725089870;
array[20675]=30'd453529185;
array[20676]=30'd473528913;
array[20677]=30'd473528913;
array[20678]=30'd473528913;
array[20679]=30'd487155275;
array[20680]=30'd473528913;
array[20681]=30'd412708426;
array[20682]=30'd460936768;
array[20683]=30'd473528913;
array[20684]=30'd487155275;
array[20685]=30'd487155275;
array[20686]=30'd487155275;
array[20687]=30'd487155275;
array[20688]=30'd487155275;
array[20689]=30'd487155275;
array[20690]=30'd473528913;
array[20691]=30'd473528913;
array[20692]=30'd412708426;
array[20693]=30'd360280652;
array[20694]=30'd460936768;
array[20695]=30'd473528913;
array[20696]=30'd360280652;
array[20697]=30'd460936768;
array[20698]=30'd473528913;
array[20699]=30'd473528913;
array[20700]=30'd473528913;
array[20701]=30'd487155275;
array[20702]=30'd487155275;
array[20703]=30'd523825734;
array[20704]=30'd697839152;
array[20705]=30'd751243845;
array[20706]=30'd792119862;
array[20707]=30'd751243845;
array[20708]=30'd483930653;
array[20709]=30'd492371499;
array[20710]=30'd492371499;
array[20711]=30'd483930653;
array[20712]=30'd804744750;
array[20713]=30'd804744750;
array[20714]=30'd804744750;
array[20715]=30'd591943231;
array[20716]=30'd483946067;
array[20717]=30'd460936768;
array[20718]=30'd473528913;
array[20719]=30'd473528913;
array[20720]=30'd473528913;
array[20721]=30'd460936768;
array[20722]=30'd412708426;
array[20723]=30'd857217603;
array[20724]=30'd959930934;
array[20725]=30'd996656669;
array[20726]=30'd916977147;
array[20727]=30'd767069629;
array[20728]=30'd876132737;
array[20729]=30'd876132737;
array[20730]=30'd766030218;
array[20731]=30'd849905057;
array[20732]=30'd945318330;
array[20733]=30'd893925805;
array[20734]=30'd778590630;
array[20735]=30'd767069629;


end

always @ (posedge clk_i) begin
	if (cen_i) begin
		val1_d1 <= array [addr_i];
		val1_d2 <= val1_d1;
		
		val2_d1 <= array2 [addr_i];
		val2_d2 <= val2_d1;
   end
end

assign val1_o = val1_d2;
assign val2_o = val2_d2;

endmodule